module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh0); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh0); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@267.2]
  input   clock, // @[:@268.4]
  input   reset, // @[:@269.4]
  input   io_enable, // @[:@270.4]
  output  io_done, // @[:@270.4]
  input   io_rst, // @[:@270.4]
  input   io_ctrDone, // @[:@270.4]
  output  io_datapathEn, // @[:@270.4]
  output  io_ctrInc // @[:@270.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@272.4]
  wire  active_reset; // @[Controllers.scala 261:22:@272.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@272.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@272.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@272.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@272.4]
  wire  done_clock; // @[Controllers.scala 262:20:@275.4]
  wire  done_reset; // @[Controllers.scala 262:20:@275.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@275.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@275.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@275.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@275.4]
  wire  RetimeWrapper_clock; // @[package.scala 98:22:@329.4]
  wire  RetimeWrapper_reset; // @[package.scala 98:22:@329.4]
  wire  RetimeWrapper_io_in; // @[package.scala 98:22:@329.4]
  wire  RetimeWrapper_io_out; // @[package.scala 98:22:@329.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 98:22:@337.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 98:22:@337.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 98:22:@337.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 98:22:@337.4]
  wire  _T_78; // @[Controllers.scala 264:38:@278.4]
  wire  _T_79; // @[Controllers.scala 264:36:@279.4]
  wire  _T_80; // @[Controllers.scala 264:48:@280.4]
  wire  _T_81; // @[Controllers.scala 264:46:@281.4]
  wire  _T_82; // @[Controllers.scala 264:62:@282.4]
  wire  _T_100; // @[package.scala 105:49:@300.4]
  reg  _T_103; // @[package.scala 53:56:@301.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 105:49:@309.4]
  wire  _T_116; // @[Controllers.scala 283:41:@317.4]
  reg  _T_125; // @[package.scala 53:56:@325.4]
  reg [31:0] _RAND_1;
  SRFF active ( // @[Controllers.scala 261:22:@272.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@275.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 98:22:@329.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 98:22:@337.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_78 = io_rst == 1'h0; // @[Controllers.scala 264:38:@278.4]
  assign _T_79 = io_enable & _T_78; // @[Controllers.scala 264:36:@279.4]
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@280.4]
  assign _T_81 = _T_79 & _T_80; // @[Controllers.scala 264:46:@281.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@282.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 105:49:@300.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 105:49:@309.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@317.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@328.4]
  assign io_datapathEn = _T_116 & io_enable; // @[Controllers.scala 283:21:@320.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@323.4]
  assign active_clock = clock; // @[:@273.4]
  assign active_reset = reset; // @[:@274.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@285.4]
  assign active_io_input_reset = io_ctrDone | io_rst; // @[Controllers.scala 265:25:@289.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@290.4]
  assign done_clock = clock; // @[:@276.4]
  assign done_reset = reset; // @[:@277.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@305.4]
  assign done_io_input_reset = io_rst; // @[Controllers.scala 267:23:@298.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@299.4]
  assign RetimeWrapper_clock = clock; // @[:@330.4]
  assign RetimeWrapper_reset = reset; // @[:@331.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 99:16:@332.4]
  assign RetimeWrapper_1_clock = clock; // @[:@338.4]
  assign RetimeWrapper_1_reset = reset; // @[:@339.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 99:16:@340.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
  end
endmodule
module fix2fixBox( // @[:@398.2]
  input  [31:0] io_a, // @[:@401.4]
  output [32:0] io_b // @[:@401.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@408.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@408.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@413.4]
endmodule
module _( // @[:@415.2]
  input  [31:0] io_b, // @[:@418.4]
  output [32:0] io_result // @[:@418.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@423.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@423.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@423.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 706:17:@431.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@426.4]
endmodule
module fix2fixBox_2( // @[:@468.2]
  input  [32:0] io_a, // @[:@471.4]
  output [31:0] io_b // @[:@471.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@481.4]
endmodule
module x38_sum( // @[:@483.2]
  input  [31:0] io_a, // @[:@486.4]
  output [31:0] io_result // @[:@486.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@494.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@494.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@501.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@501.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@519.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@519.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@499.4 Math.scala 713:14:@500.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@506.4 Math.scala 713:14:@507.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@508.4]
  _ _ ( // @[Math.scala 709:24:@494.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@501.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_2 fix2fixBox ( // @[Math.scala 141:30:@519.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@499.4 Math.scala 713:14:@500.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@506.4 Math.scala 713:14:@507.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@508.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@527.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@497.4]
  assign __1_io_b = 32'h4; // @[Math.scala 710:17:@504.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@522.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@529.2]
  input  [63:0] io_in_x32_x, // @[:@532.4]
  output        io_in_x33_y_port_0_valid, // @[:@532.4]
  output [63:0] io_in_x33_y_port_0_bits, // @[:@532.4]
  input         io_sigsIn_datapathEn // @[:@532.4]
);
  wire [31:0] x38_sum_1_io_a; // @[Math.scala 150:24:@551.4]
  wire [31:0] x38_sum_1_io_result; // @[Math.scala 150:24:@551.4]
  wire [31:0] x38_sum_number; // @[Math.scala 154:22:@557.4 Math.scala 155:14:@558.4]
  wire  _T_148; // @[FixedPoint.scala 50:25:@560.4]
  wire [31:0] _T_152; // @[Bitwise.scala 72:12:@562.4]
  x38_sum x38_sum_1 ( // @[Math.scala 150:24:@551.4]
    .io_a(x38_sum_1_io_a),
    .io_result(x38_sum_1_io_result)
  );
  assign x38_sum_number = x38_sum_1_io_result; // @[Math.scala 154:22:@557.4 Math.scala 155:14:@558.4]
  assign _T_148 = x38_sum_number[31]; // @[FixedPoint.scala 50:25:@560.4]
  assign _T_152 = _T_148 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@562.4]
  assign io_in_x33_y_port_0_valid = io_sigsIn_datapathEn; // @[MemInterfaceType.scala 311:132:@567.4]
  assign io_in_x33_y_port_0_bits = {_T_152,x38_sum_number}; // @[MemInterfaceType.scala 311:109:@566.4]
  assign x38_sum_1_io_a = io_in_x32_x[31:0]; // @[Math.scala 151:17:@554.4]
endmodule
module AccelTop( // @[:@569.2]
  input         clock, // @[:@570.4]
  input         reset, // @[:@571.4]
  input         io_enable, // @[:@572.4]
  output        io_done, // @[:@572.4]
  input  [63:0] io_argIns_0, // @[:@572.4]
  output        io_argOuts_0_port_valid, // @[:@572.4]
  output [63:0] io_argOuts_0_port_bits // @[:@572.4]
);
  wire  SingleCounter_clock; // @[Main.scala 32:32:@672.4]
  wire  SingleCounter_reset; // @[Main.scala 32:32:@672.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 32:32:@672.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 32:32:@672.4]
  wire  RetimeWrapper_clock; // @[package.scala 98:22:@690.4]
  wire  RetimeWrapper_reset; // @[package.scala 98:22:@690.4]
  wire  RetimeWrapper_io_in; // @[package.scala 98:22:@690.4]
  wire  RetimeWrapper_io_out; // @[package.scala 98:22:@690.4]
  wire  SRFF_clock; // @[Main.scala 36:28:@699.4]
  wire  SRFF_reset; // @[Main.scala 36:28:@699.4]
  wire  SRFF_io_input_set; // @[Main.scala 36:28:@699.4]
  wire  SRFF_io_input_reset; // @[Main.scala 36:28:@699.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 36:28:@699.4]
  wire  SRFF_io_output; // @[Main.scala 36:28:@699.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_datapathEn; // @[sm_RootController.scala 32:18:@737.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@737.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 98:22:@769.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 98:22:@769.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 98:22:@769.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 98:22:@769.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x32_x; // @[sm_RootController.scala 67:24:@828.4]
  wire  RootController_kernelRootController_concrete1_io_in_x33_y_port_0_valid; // @[sm_RootController.scala 67:24:@828.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x33_y_port_0_bits; // @[sm_RootController.scala 67:24:@828.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_datapathEn; // @[sm_RootController.scala 67:24:@828.4]
  wire  _T_523; // @[package.scala 101:25:@695.4 package.scala 101:25:@696.4]
  wire  _T_588; // @[Main.scala 38:44:@765.4]
  wire  _T_589; // @[Main.scala 38:53:@766.4]
  wire  _T_601; // @[package.scala 105:49:@786.4]
  reg  _T_604; // @[package.scala 53:56:@787.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 32:32:@672.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 98:22:@690.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 36:28:@699.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@737.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_datapathEn(RootController_sm_io_datapathEn),
    .io_ctrInc(RootController_sm_io_ctrInc)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 98:22:@769.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 67:24:@828.4]
    .io_in_x32_x(RootController_kernelRootController_concrete1_io_in_x32_x),
    .io_in_x33_y_port_0_valid(RootController_kernelRootController_concrete1_io_in_x33_y_port_0_valid),
    .io_in_x33_y_port_0_bits(RootController_kernelRootController_concrete1_io_in_x33_y_port_0_bits),
    .io_sigsIn_datapathEn(RootController_kernelRootController_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_523 = RetimeWrapper_io_out; // @[package.scala 101:25:@695.4 package.scala 101:25:@696.4]
  assign _T_588 = io_enable & _T_523; // @[Main.scala 38:44:@765.4]
  assign _T_589 = ~ SRFF_io_output; // @[Main.scala 38:53:@766.4]
  assign _T_601 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 105:49:@786.4]
  assign io_done = SRFF_io_output; // @[Main.scala 45:17:@785.4]
  assign io_argOuts_0_port_valid = RootController_kernelRootController_concrete1_io_in_x33_y_port_0_valid; // @[Main.scala 28:57:@668.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_x33_y_port_0_bits; // @[Main.scala 29:56:@669.4]
  assign SingleCounter_clock = clock; // @[:@673.4]
  assign SingleCounter_reset = reset; // @[:@674.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 33:79:@688.4]
  assign RetimeWrapper_clock = clock; // @[:@691.4]
  assign RetimeWrapper_reset = reset; // @[:@692.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 99:16:@693.4]
  assign SRFF_clock = clock; // @[:@700.4]
  assign SRFF_reset = reset; // @[:@701.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 54:29:@895.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 43:31:@783.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 44:36:@784.4]
  assign RootController_sm_clock = clock; // @[:@738.4]
  assign RootController_sm_reset = reset; // @[:@739.4]
  assign RootController_sm_io_enable = _T_588 & _T_589; // @[Main.scala 42:33:@782.4 SpatialBlocks.scala 112:18:@816.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@810.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_604; // @[Main.scala 46:34:@790.4]
  assign RetimeWrapper_1_clock = clock; // @[:@770.4]
  assign RetimeWrapper_1_reset = reset; // @[:@771.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 99:16:@772.4]
  assign RootController_kernelRootController_concrete1_io_in_x32_x = io_argIns_0; // @[sm_RootController.scala 48:24:@863.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_datapathEn = RootController_sm_io_datapathEn; // @[sm_RootController.scala 71:22:@881.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_604 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_604 <= 1'h0;
    end else begin
      _T_604 <= _T_601;
    end
  end
endmodule
module RetimeWrapper_4( // @[:@2605.2]
  input         clock, // @[:@2606.4]
  input         reset, // @[:@2607.4]
  input         io_flow, // @[:@2608.4]
  input  [63:0] io_in, // @[:@2608.4]
  output [63:0] io_out // @[:@2608.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2610.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@2610.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2623.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2622.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@2621.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2620.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2619.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2617.4]
endmodule
module FringeFF( // @[:@2625.2]
  input         clock, // @[:@2626.4]
  input         reset, // @[:@2627.4]
  input  [63:0] io_in, // @[:@2628.4]
  input         io_reset, // @[:@2628.4]
  output [63:0] io_out, // @[:@2628.4]
  input         io_enable // @[:@2628.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 98:22:@2631.4]
  wire  RetimeWrapper_reset; // @[package.scala 98:22:@2631.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 98:22:@2631.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 98:22:@2631.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 98:22:@2631.4]
  wire [63:0] _T_18; // @[package.scala 101:25:@2636.4 package.scala 101:25:@2637.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@2642.6]
  RetimeWrapper_4 RetimeWrapper ( // @[package.scala 98:22:@2631.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 101:25:@2636.4 package.scala 101:25:@2637.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@2642.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@2648.4]
  assign RetimeWrapper_clock = clock; // @[:@2632.4]
  assign RetimeWrapper_reset = reset; // @[:@2633.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 100:18:@2635.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 99:16:@2634.4]
endmodule
module RegFile( // @[:@31271.2]
  input         clock, // @[:@31272.4]
  input         reset, // @[:@31273.4]
  input         io_reset, // @[:@31274.4]
  output [63:0] io_argIns_0, // @[:@31274.4]
  output [63:0] io_argIns_1, // @[:@31274.4]
  output [63:0] io_argIns_2, // @[:@31274.4]
  input         io_argOuts_0_valid, // @[:@31274.4]
  input  [63:0] io_argOuts_0_bits, // @[:@31274.4]
  input         io_argOuts_1_valid, // @[:@31274.4]
  input  [63:0] io_argOuts_1_bits // @[:@31274.4]
);
  wire  regs_0_clock; // @[RegFile.scala 65:20:@33284.4]
  wire  regs_0_reset; // @[RegFile.scala 65:20:@33284.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 65:20:@33284.4]
  wire  regs_0_io_reset; // @[RegFile.scala 65:20:@33284.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 65:20:@33284.4]
  wire  regs_0_io_enable; // @[RegFile.scala 65:20:@33284.4]
  wire  regs_1_clock; // @[RegFile.scala 65:20:@33296.4]
  wire  regs_1_reset; // @[RegFile.scala 65:20:@33296.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 65:20:@33296.4]
  wire  regs_1_io_reset; // @[RegFile.scala 65:20:@33296.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 65:20:@33296.4]
  wire  regs_1_io_enable; // @[RegFile.scala 65:20:@33296.4]
  wire  regs_2_clock; // @[RegFile.scala 65:20:@33315.4]
  wire  regs_2_reset; // @[RegFile.scala 65:20:@33315.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 65:20:@33315.4]
  wire  regs_2_io_reset; // @[RegFile.scala 65:20:@33315.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 65:20:@33315.4]
  wire  regs_2_io_enable; // @[RegFile.scala 65:20:@33315.4]
  wire  regs_3_clock; // @[RegFile.scala 65:20:@33327.4]
  wire  regs_3_reset; // @[RegFile.scala 65:20:@33327.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 65:20:@33327.4]
  wire  regs_3_io_reset; // @[RegFile.scala 65:20:@33327.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 65:20:@33327.4]
  wire  regs_3_io_enable; // @[RegFile.scala 65:20:@33327.4]
  wire  regs_4_clock; // @[RegFile.scala 65:20:@33341.4]
  wire  regs_4_reset; // @[RegFile.scala 65:20:@33341.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 65:20:@33341.4]
  wire  regs_4_io_reset; // @[RegFile.scala 65:20:@33341.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 65:20:@33341.4]
  wire  regs_4_io_enable; // @[RegFile.scala 65:20:@33341.4]
  wire  regs_5_clock; // @[RegFile.scala 65:20:@33355.4]
  wire  regs_5_reset; // @[RegFile.scala 65:20:@33355.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 65:20:@33355.4]
  wire  regs_5_io_reset; // @[RegFile.scala 65:20:@33355.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 65:20:@33355.4]
  wire  regs_5_io_enable; // @[RegFile.scala 65:20:@33355.4]
  wire  regs_6_clock; // @[RegFile.scala 65:20:@33369.4]
  wire  regs_6_reset; // @[RegFile.scala 65:20:@33369.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 65:20:@33369.4]
  wire  regs_6_io_reset; // @[RegFile.scala 65:20:@33369.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 65:20:@33369.4]
  wire  regs_6_io_enable; // @[RegFile.scala 65:20:@33369.4]
  wire  regs_7_clock; // @[RegFile.scala 65:20:@33383.4]
  wire  regs_7_reset; // @[RegFile.scala 65:20:@33383.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 65:20:@33383.4]
  wire  regs_7_io_reset; // @[RegFile.scala 65:20:@33383.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 65:20:@33383.4]
  wire  regs_7_io_enable; // @[RegFile.scala 65:20:@33383.4]
  wire  regs_8_clock; // @[RegFile.scala 65:20:@33397.4]
  wire  regs_8_reset; // @[RegFile.scala 65:20:@33397.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 65:20:@33397.4]
  wire  regs_8_io_reset; // @[RegFile.scala 65:20:@33397.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 65:20:@33397.4]
  wire  regs_8_io_enable; // @[RegFile.scala 65:20:@33397.4]
  wire  regs_9_clock; // @[RegFile.scala 65:20:@33411.4]
  wire  regs_9_reset; // @[RegFile.scala 65:20:@33411.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 65:20:@33411.4]
  wire  regs_9_io_reset; // @[RegFile.scala 65:20:@33411.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 65:20:@33411.4]
  wire  regs_9_io_enable; // @[RegFile.scala 65:20:@33411.4]
  wire  regs_10_clock; // @[RegFile.scala 65:20:@33425.4]
  wire  regs_10_reset; // @[RegFile.scala 65:20:@33425.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 65:20:@33425.4]
  wire  regs_10_io_reset; // @[RegFile.scala 65:20:@33425.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 65:20:@33425.4]
  wire  regs_10_io_enable; // @[RegFile.scala 65:20:@33425.4]
  wire  regs_11_clock; // @[RegFile.scala 65:20:@33439.4]
  wire  regs_11_reset; // @[RegFile.scala 65:20:@33439.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 65:20:@33439.4]
  wire  regs_11_io_reset; // @[RegFile.scala 65:20:@33439.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 65:20:@33439.4]
  wire  regs_11_io_enable; // @[RegFile.scala 65:20:@33439.4]
  wire  regs_12_clock; // @[RegFile.scala 65:20:@33453.4]
  wire  regs_12_reset; // @[RegFile.scala 65:20:@33453.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 65:20:@33453.4]
  wire  regs_12_io_reset; // @[RegFile.scala 65:20:@33453.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 65:20:@33453.4]
  wire  regs_12_io_enable; // @[RegFile.scala 65:20:@33453.4]
  wire  regs_13_clock; // @[RegFile.scala 65:20:@33467.4]
  wire  regs_13_reset; // @[RegFile.scala 65:20:@33467.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 65:20:@33467.4]
  wire  regs_13_io_reset; // @[RegFile.scala 65:20:@33467.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 65:20:@33467.4]
  wire  regs_13_io_enable; // @[RegFile.scala 65:20:@33467.4]
  wire  regs_14_clock; // @[RegFile.scala 65:20:@33481.4]
  wire  regs_14_reset; // @[RegFile.scala 65:20:@33481.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 65:20:@33481.4]
  wire  regs_14_io_reset; // @[RegFile.scala 65:20:@33481.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 65:20:@33481.4]
  wire  regs_14_io_enable; // @[RegFile.scala 65:20:@33481.4]
  wire  regs_15_clock; // @[RegFile.scala 65:20:@33495.4]
  wire  regs_15_reset; // @[RegFile.scala 65:20:@33495.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 65:20:@33495.4]
  wire  regs_15_io_reset; // @[RegFile.scala 65:20:@33495.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 65:20:@33495.4]
  wire  regs_15_io_enable; // @[RegFile.scala 65:20:@33495.4]
  wire  regs_16_clock; // @[RegFile.scala 65:20:@33509.4]
  wire  regs_16_reset; // @[RegFile.scala 65:20:@33509.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 65:20:@33509.4]
  wire  regs_16_io_reset; // @[RegFile.scala 65:20:@33509.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 65:20:@33509.4]
  wire  regs_16_io_enable; // @[RegFile.scala 65:20:@33509.4]
  wire  regs_17_clock; // @[RegFile.scala 65:20:@33523.4]
  wire  regs_17_reset; // @[RegFile.scala 65:20:@33523.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 65:20:@33523.4]
  wire  regs_17_io_reset; // @[RegFile.scala 65:20:@33523.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 65:20:@33523.4]
  wire  regs_17_io_enable; // @[RegFile.scala 65:20:@33523.4]
  wire  regs_18_clock; // @[RegFile.scala 65:20:@33537.4]
  wire  regs_18_reset; // @[RegFile.scala 65:20:@33537.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 65:20:@33537.4]
  wire  regs_18_io_reset; // @[RegFile.scala 65:20:@33537.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 65:20:@33537.4]
  wire  regs_18_io_enable; // @[RegFile.scala 65:20:@33537.4]
  wire  regs_19_clock; // @[RegFile.scala 65:20:@33551.4]
  wire  regs_19_reset; // @[RegFile.scala 65:20:@33551.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 65:20:@33551.4]
  wire  regs_19_io_reset; // @[RegFile.scala 65:20:@33551.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 65:20:@33551.4]
  wire  regs_19_io_enable; // @[RegFile.scala 65:20:@33551.4]
  wire  regs_20_clock; // @[RegFile.scala 65:20:@33565.4]
  wire  regs_20_reset; // @[RegFile.scala 65:20:@33565.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 65:20:@33565.4]
  wire  regs_20_io_reset; // @[RegFile.scala 65:20:@33565.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 65:20:@33565.4]
  wire  regs_20_io_enable; // @[RegFile.scala 65:20:@33565.4]
  wire  regs_21_clock; // @[RegFile.scala 65:20:@33579.4]
  wire  regs_21_reset; // @[RegFile.scala 65:20:@33579.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 65:20:@33579.4]
  wire  regs_21_io_reset; // @[RegFile.scala 65:20:@33579.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 65:20:@33579.4]
  wire  regs_21_io_enable; // @[RegFile.scala 65:20:@33579.4]
  wire  regs_22_clock; // @[RegFile.scala 65:20:@33593.4]
  wire  regs_22_reset; // @[RegFile.scala 65:20:@33593.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 65:20:@33593.4]
  wire  regs_22_io_reset; // @[RegFile.scala 65:20:@33593.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 65:20:@33593.4]
  wire  regs_22_io_enable; // @[RegFile.scala 65:20:@33593.4]
  wire  regs_23_clock; // @[RegFile.scala 65:20:@33607.4]
  wire  regs_23_reset; // @[RegFile.scala 65:20:@33607.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 65:20:@33607.4]
  wire  regs_23_io_reset; // @[RegFile.scala 65:20:@33607.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 65:20:@33607.4]
  wire  regs_23_io_enable; // @[RegFile.scala 65:20:@33607.4]
  wire  regs_24_clock; // @[RegFile.scala 65:20:@33621.4]
  wire  regs_24_reset; // @[RegFile.scala 65:20:@33621.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 65:20:@33621.4]
  wire  regs_24_io_reset; // @[RegFile.scala 65:20:@33621.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 65:20:@33621.4]
  wire  regs_24_io_enable; // @[RegFile.scala 65:20:@33621.4]
  wire  regs_25_clock; // @[RegFile.scala 65:20:@33635.4]
  wire  regs_25_reset; // @[RegFile.scala 65:20:@33635.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 65:20:@33635.4]
  wire  regs_25_io_reset; // @[RegFile.scala 65:20:@33635.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 65:20:@33635.4]
  wire  regs_25_io_enable; // @[RegFile.scala 65:20:@33635.4]
  wire  regs_26_clock; // @[RegFile.scala 65:20:@33649.4]
  wire  regs_26_reset; // @[RegFile.scala 65:20:@33649.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 65:20:@33649.4]
  wire  regs_26_io_reset; // @[RegFile.scala 65:20:@33649.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 65:20:@33649.4]
  wire  regs_26_io_enable; // @[RegFile.scala 65:20:@33649.4]
  wire  regs_27_clock; // @[RegFile.scala 65:20:@33663.4]
  wire  regs_27_reset; // @[RegFile.scala 65:20:@33663.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 65:20:@33663.4]
  wire  regs_27_io_reset; // @[RegFile.scala 65:20:@33663.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 65:20:@33663.4]
  wire  regs_27_io_enable; // @[RegFile.scala 65:20:@33663.4]
  wire  regs_28_clock; // @[RegFile.scala 65:20:@33677.4]
  wire  regs_28_reset; // @[RegFile.scala 65:20:@33677.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 65:20:@33677.4]
  wire  regs_28_io_reset; // @[RegFile.scala 65:20:@33677.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 65:20:@33677.4]
  wire  regs_28_io_enable; // @[RegFile.scala 65:20:@33677.4]
  wire  regs_29_clock; // @[RegFile.scala 65:20:@33691.4]
  wire  regs_29_reset; // @[RegFile.scala 65:20:@33691.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 65:20:@33691.4]
  wire  regs_29_io_reset; // @[RegFile.scala 65:20:@33691.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 65:20:@33691.4]
  wire  regs_29_io_enable; // @[RegFile.scala 65:20:@33691.4]
  wire  regs_30_clock; // @[RegFile.scala 65:20:@33705.4]
  wire  regs_30_reset; // @[RegFile.scala 65:20:@33705.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 65:20:@33705.4]
  wire  regs_30_io_reset; // @[RegFile.scala 65:20:@33705.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 65:20:@33705.4]
  wire  regs_30_io_enable; // @[RegFile.scala 65:20:@33705.4]
  wire  regs_31_clock; // @[RegFile.scala 65:20:@33719.4]
  wire  regs_31_reset; // @[RegFile.scala 65:20:@33719.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 65:20:@33719.4]
  wire  regs_31_io_reset; // @[RegFile.scala 65:20:@33719.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 65:20:@33719.4]
  wire  regs_31_io_enable; // @[RegFile.scala 65:20:@33719.4]
  wire  regs_32_clock; // @[RegFile.scala 65:20:@33733.4]
  wire  regs_32_reset; // @[RegFile.scala 65:20:@33733.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 65:20:@33733.4]
  wire  regs_32_io_reset; // @[RegFile.scala 65:20:@33733.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 65:20:@33733.4]
  wire  regs_32_io_enable; // @[RegFile.scala 65:20:@33733.4]
  wire  regs_33_clock; // @[RegFile.scala 65:20:@33747.4]
  wire  regs_33_reset; // @[RegFile.scala 65:20:@33747.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 65:20:@33747.4]
  wire  regs_33_io_reset; // @[RegFile.scala 65:20:@33747.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 65:20:@33747.4]
  wire  regs_33_io_enable; // @[RegFile.scala 65:20:@33747.4]
  wire  regs_34_clock; // @[RegFile.scala 65:20:@33761.4]
  wire  regs_34_reset; // @[RegFile.scala 65:20:@33761.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 65:20:@33761.4]
  wire  regs_34_io_reset; // @[RegFile.scala 65:20:@33761.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 65:20:@33761.4]
  wire  regs_34_io_enable; // @[RegFile.scala 65:20:@33761.4]
  wire  regs_35_clock; // @[RegFile.scala 65:20:@33775.4]
  wire  regs_35_reset; // @[RegFile.scala 65:20:@33775.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 65:20:@33775.4]
  wire  regs_35_io_reset; // @[RegFile.scala 65:20:@33775.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 65:20:@33775.4]
  wire  regs_35_io_enable; // @[RegFile.scala 65:20:@33775.4]
  wire  regs_36_clock; // @[RegFile.scala 65:20:@33789.4]
  wire  regs_36_reset; // @[RegFile.scala 65:20:@33789.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 65:20:@33789.4]
  wire  regs_36_io_reset; // @[RegFile.scala 65:20:@33789.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 65:20:@33789.4]
  wire  regs_36_io_enable; // @[RegFile.scala 65:20:@33789.4]
  wire  regs_37_clock; // @[RegFile.scala 65:20:@33803.4]
  wire  regs_37_reset; // @[RegFile.scala 65:20:@33803.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 65:20:@33803.4]
  wire  regs_37_io_reset; // @[RegFile.scala 65:20:@33803.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 65:20:@33803.4]
  wire  regs_37_io_enable; // @[RegFile.scala 65:20:@33803.4]
  wire  regs_38_clock; // @[RegFile.scala 65:20:@33817.4]
  wire  regs_38_reset; // @[RegFile.scala 65:20:@33817.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 65:20:@33817.4]
  wire  regs_38_io_reset; // @[RegFile.scala 65:20:@33817.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 65:20:@33817.4]
  wire  regs_38_io_enable; // @[RegFile.scala 65:20:@33817.4]
  wire  regs_39_clock; // @[RegFile.scala 65:20:@33831.4]
  wire  regs_39_reset; // @[RegFile.scala 65:20:@33831.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 65:20:@33831.4]
  wire  regs_39_io_reset; // @[RegFile.scala 65:20:@33831.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 65:20:@33831.4]
  wire  regs_39_io_enable; // @[RegFile.scala 65:20:@33831.4]
  wire  regs_40_clock; // @[RegFile.scala 65:20:@33845.4]
  wire  regs_40_reset; // @[RegFile.scala 65:20:@33845.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 65:20:@33845.4]
  wire  regs_40_io_reset; // @[RegFile.scala 65:20:@33845.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 65:20:@33845.4]
  wire  regs_40_io_enable; // @[RegFile.scala 65:20:@33845.4]
  wire  regs_41_clock; // @[RegFile.scala 65:20:@33859.4]
  wire  regs_41_reset; // @[RegFile.scala 65:20:@33859.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 65:20:@33859.4]
  wire  regs_41_io_reset; // @[RegFile.scala 65:20:@33859.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 65:20:@33859.4]
  wire  regs_41_io_enable; // @[RegFile.scala 65:20:@33859.4]
  wire  regs_42_clock; // @[RegFile.scala 65:20:@33873.4]
  wire  regs_42_reset; // @[RegFile.scala 65:20:@33873.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 65:20:@33873.4]
  wire  regs_42_io_reset; // @[RegFile.scala 65:20:@33873.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 65:20:@33873.4]
  wire  regs_42_io_enable; // @[RegFile.scala 65:20:@33873.4]
  wire  regs_43_clock; // @[RegFile.scala 65:20:@33887.4]
  wire  regs_43_reset; // @[RegFile.scala 65:20:@33887.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 65:20:@33887.4]
  wire  regs_43_io_reset; // @[RegFile.scala 65:20:@33887.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 65:20:@33887.4]
  wire  regs_43_io_enable; // @[RegFile.scala 65:20:@33887.4]
  wire  regs_44_clock; // @[RegFile.scala 65:20:@33901.4]
  wire  regs_44_reset; // @[RegFile.scala 65:20:@33901.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 65:20:@33901.4]
  wire  regs_44_io_reset; // @[RegFile.scala 65:20:@33901.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 65:20:@33901.4]
  wire  regs_44_io_enable; // @[RegFile.scala 65:20:@33901.4]
  wire  regs_45_clock; // @[RegFile.scala 65:20:@33915.4]
  wire  regs_45_reset; // @[RegFile.scala 65:20:@33915.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 65:20:@33915.4]
  wire  regs_45_io_reset; // @[RegFile.scala 65:20:@33915.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 65:20:@33915.4]
  wire  regs_45_io_enable; // @[RegFile.scala 65:20:@33915.4]
  wire  regs_46_clock; // @[RegFile.scala 65:20:@33929.4]
  wire  regs_46_reset; // @[RegFile.scala 65:20:@33929.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 65:20:@33929.4]
  wire  regs_46_io_reset; // @[RegFile.scala 65:20:@33929.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 65:20:@33929.4]
  wire  regs_46_io_enable; // @[RegFile.scala 65:20:@33929.4]
  wire  regs_47_clock; // @[RegFile.scala 65:20:@33943.4]
  wire  regs_47_reset; // @[RegFile.scala 65:20:@33943.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 65:20:@33943.4]
  wire  regs_47_io_reset; // @[RegFile.scala 65:20:@33943.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 65:20:@33943.4]
  wire  regs_47_io_enable; // @[RegFile.scala 65:20:@33943.4]
  wire  regs_48_clock; // @[RegFile.scala 65:20:@33957.4]
  wire  regs_48_reset; // @[RegFile.scala 65:20:@33957.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 65:20:@33957.4]
  wire  regs_48_io_reset; // @[RegFile.scala 65:20:@33957.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 65:20:@33957.4]
  wire  regs_48_io_enable; // @[RegFile.scala 65:20:@33957.4]
  wire  regs_49_clock; // @[RegFile.scala 65:20:@33971.4]
  wire  regs_49_reset; // @[RegFile.scala 65:20:@33971.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 65:20:@33971.4]
  wire  regs_49_io_reset; // @[RegFile.scala 65:20:@33971.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 65:20:@33971.4]
  wire  regs_49_io_enable; // @[RegFile.scala 65:20:@33971.4]
  wire  regs_50_clock; // @[RegFile.scala 65:20:@33985.4]
  wire  regs_50_reset; // @[RegFile.scala 65:20:@33985.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 65:20:@33985.4]
  wire  regs_50_io_reset; // @[RegFile.scala 65:20:@33985.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 65:20:@33985.4]
  wire  regs_50_io_enable; // @[RegFile.scala 65:20:@33985.4]
  wire  regs_51_clock; // @[RegFile.scala 65:20:@33999.4]
  wire  regs_51_reset; // @[RegFile.scala 65:20:@33999.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 65:20:@33999.4]
  wire  regs_51_io_reset; // @[RegFile.scala 65:20:@33999.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 65:20:@33999.4]
  wire  regs_51_io_enable; // @[RegFile.scala 65:20:@33999.4]
  wire  regs_52_clock; // @[RegFile.scala 65:20:@34013.4]
  wire  regs_52_reset; // @[RegFile.scala 65:20:@34013.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 65:20:@34013.4]
  wire  regs_52_io_reset; // @[RegFile.scala 65:20:@34013.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 65:20:@34013.4]
  wire  regs_52_io_enable; // @[RegFile.scala 65:20:@34013.4]
  wire  regs_53_clock; // @[RegFile.scala 65:20:@34027.4]
  wire  regs_53_reset; // @[RegFile.scala 65:20:@34027.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 65:20:@34027.4]
  wire  regs_53_io_reset; // @[RegFile.scala 65:20:@34027.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 65:20:@34027.4]
  wire  regs_53_io_enable; // @[RegFile.scala 65:20:@34027.4]
  wire  regs_54_clock; // @[RegFile.scala 65:20:@34041.4]
  wire  regs_54_reset; // @[RegFile.scala 65:20:@34041.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 65:20:@34041.4]
  wire  regs_54_io_reset; // @[RegFile.scala 65:20:@34041.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 65:20:@34041.4]
  wire  regs_54_io_enable; // @[RegFile.scala 65:20:@34041.4]
  wire  regs_55_clock; // @[RegFile.scala 65:20:@34055.4]
  wire  regs_55_reset; // @[RegFile.scala 65:20:@34055.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 65:20:@34055.4]
  wire  regs_55_io_reset; // @[RegFile.scala 65:20:@34055.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 65:20:@34055.4]
  wire  regs_55_io_enable; // @[RegFile.scala 65:20:@34055.4]
  wire  regs_56_clock; // @[RegFile.scala 65:20:@34069.4]
  wire  regs_56_reset; // @[RegFile.scala 65:20:@34069.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 65:20:@34069.4]
  wire  regs_56_io_reset; // @[RegFile.scala 65:20:@34069.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 65:20:@34069.4]
  wire  regs_56_io_enable; // @[RegFile.scala 65:20:@34069.4]
  wire  regs_57_clock; // @[RegFile.scala 65:20:@34083.4]
  wire  regs_57_reset; // @[RegFile.scala 65:20:@34083.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 65:20:@34083.4]
  wire  regs_57_io_reset; // @[RegFile.scala 65:20:@34083.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 65:20:@34083.4]
  wire  regs_57_io_enable; // @[RegFile.scala 65:20:@34083.4]
  wire  regs_58_clock; // @[RegFile.scala 65:20:@34097.4]
  wire  regs_58_reset; // @[RegFile.scala 65:20:@34097.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 65:20:@34097.4]
  wire  regs_58_io_reset; // @[RegFile.scala 65:20:@34097.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 65:20:@34097.4]
  wire  regs_58_io_enable; // @[RegFile.scala 65:20:@34097.4]
  wire  regs_59_clock; // @[RegFile.scala 65:20:@34111.4]
  wire  regs_59_reset; // @[RegFile.scala 65:20:@34111.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 65:20:@34111.4]
  wire  regs_59_io_reset; // @[RegFile.scala 65:20:@34111.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 65:20:@34111.4]
  wire  regs_59_io_enable; // @[RegFile.scala 65:20:@34111.4]
  wire  regs_60_clock; // @[RegFile.scala 65:20:@34125.4]
  wire  regs_60_reset; // @[RegFile.scala 65:20:@34125.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 65:20:@34125.4]
  wire  regs_60_io_reset; // @[RegFile.scala 65:20:@34125.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 65:20:@34125.4]
  wire  regs_60_io_enable; // @[RegFile.scala 65:20:@34125.4]
  wire  regs_61_clock; // @[RegFile.scala 65:20:@34139.4]
  wire  regs_61_reset; // @[RegFile.scala 65:20:@34139.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 65:20:@34139.4]
  wire  regs_61_io_reset; // @[RegFile.scala 65:20:@34139.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 65:20:@34139.4]
  wire  regs_61_io_enable; // @[RegFile.scala 65:20:@34139.4]
  wire  regs_62_clock; // @[RegFile.scala 65:20:@34153.4]
  wire  regs_62_reset; // @[RegFile.scala 65:20:@34153.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 65:20:@34153.4]
  wire  regs_62_io_reset; // @[RegFile.scala 65:20:@34153.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 65:20:@34153.4]
  wire  regs_62_io_enable; // @[RegFile.scala 65:20:@34153.4]
  wire  regs_63_clock; // @[RegFile.scala 65:20:@34167.4]
  wire  regs_63_reset; // @[RegFile.scala 65:20:@34167.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 65:20:@34167.4]
  wire  regs_63_io_reset; // @[RegFile.scala 65:20:@34167.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 65:20:@34167.4]
  wire  regs_63_io_enable; // @[RegFile.scala 65:20:@34167.4]
  wire  regs_64_clock; // @[RegFile.scala 65:20:@34181.4]
  wire  regs_64_reset; // @[RegFile.scala 65:20:@34181.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 65:20:@34181.4]
  wire  regs_64_io_reset; // @[RegFile.scala 65:20:@34181.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 65:20:@34181.4]
  wire  regs_64_io_enable; // @[RegFile.scala 65:20:@34181.4]
  wire  regs_65_clock; // @[RegFile.scala 65:20:@34195.4]
  wire  regs_65_reset; // @[RegFile.scala 65:20:@34195.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 65:20:@34195.4]
  wire  regs_65_io_reset; // @[RegFile.scala 65:20:@34195.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 65:20:@34195.4]
  wire  regs_65_io_enable; // @[RegFile.scala 65:20:@34195.4]
  wire  regs_66_clock; // @[RegFile.scala 65:20:@34209.4]
  wire  regs_66_reset; // @[RegFile.scala 65:20:@34209.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 65:20:@34209.4]
  wire  regs_66_io_reset; // @[RegFile.scala 65:20:@34209.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 65:20:@34209.4]
  wire  regs_66_io_enable; // @[RegFile.scala 65:20:@34209.4]
  wire  regs_67_clock; // @[RegFile.scala 65:20:@34223.4]
  wire  regs_67_reset; // @[RegFile.scala 65:20:@34223.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 65:20:@34223.4]
  wire  regs_67_io_reset; // @[RegFile.scala 65:20:@34223.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 65:20:@34223.4]
  wire  regs_67_io_enable; // @[RegFile.scala 65:20:@34223.4]
  wire  regs_68_clock; // @[RegFile.scala 65:20:@34237.4]
  wire  regs_68_reset; // @[RegFile.scala 65:20:@34237.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 65:20:@34237.4]
  wire  regs_68_io_reset; // @[RegFile.scala 65:20:@34237.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 65:20:@34237.4]
  wire  regs_68_io_enable; // @[RegFile.scala 65:20:@34237.4]
  wire  regs_69_clock; // @[RegFile.scala 65:20:@34251.4]
  wire  regs_69_reset; // @[RegFile.scala 65:20:@34251.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 65:20:@34251.4]
  wire  regs_69_io_reset; // @[RegFile.scala 65:20:@34251.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 65:20:@34251.4]
  wire  regs_69_io_enable; // @[RegFile.scala 65:20:@34251.4]
  wire  regs_70_clock; // @[RegFile.scala 65:20:@34265.4]
  wire  regs_70_reset; // @[RegFile.scala 65:20:@34265.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 65:20:@34265.4]
  wire  regs_70_io_reset; // @[RegFile.scala 65:20:@34265.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 65:20:@34265.4]
  wire  regs_70_io_enable; // @[RegFile.scala 65:20:@34265.4]
  wire  regs_71_clock; // @[RegFile.scala 65:20:@34279.4]
  wire  regs_71_reset; // @[RegFile.scala 65:20:@34279.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 65:20:@34279.4]
  wire  regs_71_io_reset; // @[RegFile.scala 65:20:@34279.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 65:20:@34279.4]
  wire  regs_71_io_enable; // @[RegFile.scala 65:20:@34279.4]
  wire  regs_72_clock; // @[RegFile.scala 65:20:@34293.4]
  wire  regs_72_reset; // @[RegFile.scala 65:20:@34293.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 65:20:@34293.4]
  wire  regs_72_io_reset; // @[RegFile.scala 65:20:@34293.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 65:20:@34293.4]
  wire  regs_72_io_enable; // @[RegFile.scala 65:20:@34293.4]
  wire  regs_73_clock; // @[RegFile.scala 65:20:@34307.4]
  wire  regs_73_reset; // @[RegFile.scala 65:20:@34307.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 65:20:@34307.4]
  wire  regs_73_io_reset; // @[RegFile.scala 65:20:@34307.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 65:20:@34307.4]
  wire  regs_73_io_enable; // @[RegFile.scala 65:20:@34307.4]
  wire  regs_74_clock; // @[RegFile.scala 65:20:@34321.4]
  wire  regs_74_reset; // @[RegFile.scala 65:20:@34321.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 65:20:@34321.4]
  wire  regs_74_io_reset; // @[RegFile.scala 65:20:@34321.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 65:20:@34321.4]
  wire  regs_74_io_enable; // @[RegFile.scala 65:20:@34321.4]
  wire  regs_75_clock; // @[RegFile.scala 65:20:@34335.4]
  wire  regs_75_reset; // @[RegFile.scala 65:20:@34335.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 65:20:@34335.4]
  wire  regs_75_io_reset; // @[RegFile.scala 65:20:@34335.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 65:20:@34335.4]
  wire  regs_75_io_enable; // @[RegFile.scala 65:20:@34335.4]
  wire  regs_76_clock; // @[RegFile.scala 65:20:@34349.4]
  wire  regs_76_reset; // @[RegFile.scala 65:20:@34349.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 65:20:@34349.4]
  wire  regs_76_io_reset; // @[RegFile.scala 65:20:@34349.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 65:20:@34349.4]
  wire  regs_76_io_enable; // @[RegFile.scala 65:20:@34349.4]
  wire  regs_77_clock; // @[RegFile.scala 65:20:@34363.4]
  wire  regs_77_reset; // @[RegFile.scala 65:20:@34363.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 65:20:@34363.4]
  wire  regs_77_io_reset; // @[RegFile.scala 65:20:@34363.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 65:20:@34363.4]
  wire  regs_77_io_enable; // @[RegFile.scala 65:20:@34363.4]
  wire  regs_78_clock; // @[RegFile.scala 65:20:@34377.4]
  wire  regs_78_reset; // @[RegFile.scala 65:20:@34377.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 65:20:@34377.4]
  wire  regs_78_io_reset; // @[RegFile.scala 65:20:@34377.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 65:20:@34377.4]
  wire  regs_78_io_enable; // @[RegFile.scala 65:20:@34377.4]
  wire  regs_79_clock; // @[RegFile.scala 65:20:@34391.4]
  wire  regs_79_reset; // @[RegFile.scala 65:20:@34391.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 65:20:@34391.4]
  wire  regs_79_io_reset; // @[RegFile.scala 65:20:@34391.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 65:20:@34391.4]
  wire  regs_79_io_enable; // @[RegFile.scala 65:20:@34391.4]
  wire  regs_80_clock; // @[RegFile.scala 65:20:@34405.4]
  wire  regs_80_reset; // @[RegFile.scala 65:20:@34405.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 65:20:@34405.4]
  wire  regs_80_io_reset; // @[RegFile.scala 65:20:@34405.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 65:20:@34405.4]
  wire  regs_80_io_enable; // @[RegFile.scala 65:20:@34405.4]
  wire  regs_81_clock; // @[RegFile.scala 65:20:@34419.4]
  wire  regs_81_reset; // @[RegFile.scala 65:20:@34419.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 65:20:@34419.4]
  wire  regs_81_io_reset; // @[RegFile.scala 65:20:@34419.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 65:20:@34419.4]
  wire  regs_81_io_enable; // @[RegFile.scala 65:20:@34419.4]
  wire  regs_82_clock; // @[RegFile.scala 65:20:@34433.4]
  wire  regs_82_reset; // @[RegFile.scala 65:20:@34433.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 65:20:@34433.4]
  wire  regs_82_io_reset; // @[RegFile.scala 65:20:@34433.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 65:20:@34433.4]
  wire  regs_82_io_enable; // @[RegFile.scala 65:20:@34433.4]
  wire  regs_83_clock; // @[RegFile.scala 65:20:@34447.4]
  wire  regs_83_reset; // @[RegFile.scala 65:20:@34447.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 65:20:@34447.4]
  wire  regs_83_io_reset; // @[RegFile.scala 65:20:@34447.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 65:20:@34447.4]
  wire  regs_83_io_enable; // @[RegFile.scala 65:20:@34447.4]
  wire  regs_84_clock; // @[RegFile.scala 65:20:@34461.4]
  wire  regs_84_reset; // @[RegFile.scala 65:20:@34461.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 65:20:@34461.4]
  wire  regs_84_io_reset; // @[RegFile.scala 65:20:@34461.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 65:20:@34461.4]
  wire  regs_84_io_enable; // @[RegFile.scala 65:20:@34461.4]
  wire  regs_85_clock; // @[RegFile.scala 65:20:@34475.4]
  wire  regs_85_reset; // @[RegFile.scala 65:20:@34475.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 65:20:@34475.4]
  wire  regs_85_io_reset; // @[RegFile.scala 65:20:@34475.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 65:20:@34475.4]
  wire  regs_85_io_enable; // @[RegFile.scala 65:20:@34475.4]
  wire  regs_86_clock; // @[RegFile.scala 65:20:@34489.4]
  wire  regs_86_reset; // @[RegFile.scala 65:20:@34489.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 65:20:@34489.4]
  wire  regs_86_io_reset; // @[RegFile.scala 65:20:@34489.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 65:20:@34489.4]
  wire  regs_86_io_enable; // @[RegFile.scala 65:20:@34489.4]
  wire  regs_87_clock; // @[RegFile.scala 65:20:@34503.4]
  wire  regs_87_reset; // @[RegFile.scala 65:20:@34503.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 65:20:@34503.4]
  wire  regs_87_io_reset; // @[RegFile.scala 65:20:@34503.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 65:20:@34503.4]
  wire  regs_87_io_enable; // @[RegFile.scala 65:20:@34503.4]
  wire  regs_88_clock; // @[RegFile.scala 65:20:@34517.4]
  wire  regs_88_reset; // @[RegFile.scala 65:20:@34517.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 65:20:@34517.4]
  wire  regs_88_io_reset; // @[RegFile.scala 65:20:@34517.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 65:20:@34517.4]
  wire  regs_88_io_enable; // @[RegFile.scala 65:20:@34517.4]
  wire  regs_89_clock; // @[RegFile.scala 65:20:@34531.4]
  wire  regs_89_reset; // @[RegFile.scala 65:20:@34531.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 65:20:@34531.4]
  wire  regs_89_io_reset; // @[RegFile.scala 65:20:@34531.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 65:20:@34531.4]
  wire  regs_89_io_enable; // @[RegFile.scala 65:20:@34531.4]
  wire  regs_90_clock; // @[RegFile.scala 65:20:@34545.4]
  wire  regs_90_reset; // @[RegFile.scala 65:20:@34545.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 65:20:@34545.4]
  wire  regs_90_io_reset; // @[RegFile.scala 65:20:@34545.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 65:20:@34545.4]
  wire  regs_90_io_enable; // @[RegFile.scala 65:20:@34545.4]
  wire  regs_91_clock; // @[RegFile.scala 65:20:@34559.4]
  wire  regs_91_reset; // @[RegFile.scala 65:20:@34559.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 65:20:@34559.4]
  wire  regs_91_io_reset; // @[RegFile.scala 65:20:@34559.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 65:20:@34559.4]
  wire  regs_91_io_enable; // @[RegFile.scala 65:20:@34559.4]
  wire  regs_92_clock; // @[RegFile.scala 65:20:@34573.4]
  wire  regs_92_reset; // @[RegFile.scala 65:20:@34573.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 65:20:@34573.4]
  wire  regs_92_io_reset; // @[RegFile.scala 65:20:@34573.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 65:20:@34573.4]
  wire  regs_92_io_enable; // @[RegFile.scala 65:20:@34573.4]
  wire  regs_93_clock; // @[RegFile.scala 65:20:@34587.4]
  wire  regs_93_reset; // @[RegFile.scala 65:20:@34587.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 65:20:@34587.4]
  wire  regs_93_io_reset; // @[RegFile.scala 65:20:@34587.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 65:20:@34587.4]
  wire  regs_93_io_enable; // @[RegFile.scala 65:20:@34587.4]
  wire  regs_94_clock; // @[RegFile.scala 65:20:@34601.4]
  wire  regs_94_reset; // @[RegFile.scala 65:20:@34601.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 65:20:@34601.4]
  wire  regs_94_io_reset; // @[RegFile.scala 65:20:@34601.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 65:20:@34601.4]
  wire  regs_94_io_enable; // @[RegFile.scala 65:20:@34601.4]
  wire  regs_95_clock; // @[RegFile.scala 65:20:@34615.4]
  wire  regs_95_reset; // @[RegFile.scala 65:20:@34615.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 65:20:@34615.4]
  wire  regs_95_io_reset; // @[RegFile.scala 65:20:@34615.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 65:20:@34615.4]
  wire  regs_95_io_enable; // @[RegFile.scala 65:20:@34615.4]
  wire  regs_96_clock; // @[RegFile.scala 65:20:@34629.4]
  wire  regs_96_reset; // @[RegFile.scala 65:20:@34629.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 65:20:@34629.4]
  wire  regs_96_io_reset; // @[RegFile.scala 65:20:@34629.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 65:20:@34629.4]
  wire  regs_96_io_enable; // @[RegFile.scala 65:20:@34629.4]
  wire  regs_97_clock; // @[RegFile.scala 65:20:@34643.4]
  wire  regs_97_reset; // @[RegFile.scala 65:20:@34643.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 65:20:@34643.4]
  wire  regs_97_io_reset; // @[RegFile.scala 65:20:@34643.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 65:20:@34643.4]
  wire  regs_97_io_enable; // @[RegFile.scala 65:20:@34643.4]
  wire  regs_98_clock; // @[RegFile.scala 65:20:@34657.4]
  wire  regs_98_reset; // @[RegFile.scala 65:20:@34657.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 65:20:@34657.4]
  wire  regs_98_io_reset; // @[RegFile.scala 65:20:@34657.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 65:20:@34657.4]
  wire  regs_98_io_enable; // @[RegFile.scala 65:20:@34657.4]
  wire  regs_99_clock; // @[RegFile.scala 65:20:@34671.4]
  wire  regs_99_reset; // @[RegFile.scala 65:20:@34671.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 65:20:@34671.4]
  wire  regs_99_io_reset; // @[RegFile.scala 65:20:@34671.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 65:20:@34671.4]
  wire  regs_99_io_enable; // @[RegFile.scala 65:20:@34671.4]
  wire  regs_100_clock; // @[RegFile.scala 65:20:@34685.4]
  wire  regs_100_reset; // @[RegFile.scala 65:20:@34685.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 65:20:@34685.4]
  wire  regs_100_io_reset; // @[RegFile.scala 65:20:@34685.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 65:20:@34685.4]
  wire  regs_100_io_enable; // @[RegFile.scala 65:20:@34685.4]
  wire  regs_101_clock; // @[RegFile.scala 65:20:@34699.4]
  wire  regs_101_reset; // @[RegFile.scala 65:20:@34699.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 65:20:@34699.4]
  wire  regs_101_io_reset; // @[RegFile.scala 65:20:@34699.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 65:20:@34699.4]
  wire  regs_101_io_enable; // @[RegFile.scala 65:20:@34699.4]
  wire  regs_102_clock; // @[RegFile.scala 65:20:@34713.4]
  wire  regs_102_reset; // @[RegFile.scala 65:20:@34713.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 65:20:@34713.4]
  wire  regs_102_io_reset; // @[RegFile.scala 65:20:@34713.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 65:20:@34713.4]
  wire  regs_102_io_enable; // @[RegFile.scala 65:20:@34713.4]
  wire  regs_103_clock; // @[RegFile.scala 65:20:@34727.4]
  wire  regs_103_reset; // @[RegFile.scala 65:20:@34727.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 65:20:@34727.4]
  wire  regs_103_io_reset; // @[RegFile.scala 65:20:@34727.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 65:20:@34727.4]
  wire  regs_103_io_enable; // @[RegFile.scala 65:20:@34727.4]
  wire  regs_104_clock; // @[RegFile.scala 65:20:@34741.4]
  wire  regs_104_reset; // @[RegFile.scala 65:20:@34741.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 65:20:@34741.4]
  wire  regs_104_io_reset; // @[RegFile.scala 65:20:@34741.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 65:20:@34741.4]
  wire  regs_104_io_enable; // @[RegFile.scala 65:20:@34741.4]
  wire  regs_105_clock; // @[RegFile.scala 65:20:@34755.4]
  wire  regs_105_reset; // @[RegFile.scala 65:20:@34755.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 65:20:@34755.4]
  wire  regs_105_io_reset; // @[RegFile.scala 65:20:@34755.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 65:20:@34755.4]
  wire  regs_105_io_enable; // @[RegFile.scala 65:20:@34755.4]
  wire  regs_106_clock; // @[RegFile.scala 65:20:@34769.4]
  wire  regs_106_reset; // @[RegFile.scala 65:20:@34769.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 65:20:@34769.4]
  wire  regs_106_io_reset; // @[RegFile.scala 65:20:@34769.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 65:20:@34769.4]
  wire  regs_106_io_enable; // @[RegFile.scala 65:20:@34769.4]
  wire  regs_107_clock; // @[RegFile.scala 65:20:@34783.4]
  wire  regs_107_reset; // @[RegFile.scala 65:20:@34783.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 65:20:@34783.4]
  wire  regs_107_io_reset; // @[RegFile.scala 65:20:@34783.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 65:20:@34783.4]
  wire  regs_107_io_enable; // @[RegFile.scala 65:20:@34783.4]
  wire  regs_108_clock; // @[RegFile.scala 65:20:@34797.4]
  wire  regs_108_reset; // @[RegFile.scala 65:20:@34797.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 65:20:@34797.4]
  wire  regs_108_io_reset; // @[RegFile.scala 65:20:@34797.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 65:20:@34797.4]
  wire  regs_108_io_enable; // @[RegFile.scala 65:20:@34797.4]
  wire  regs_109_clock; // @[RegFile.scala 65:20:@34811.4]
  wire  regs_109_reset; // @[RegFile.scala 65:20:@34811.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 65:20:@34811.4]
  wire  regs_109_io_reset; // @[RegFile.scala 65:20:@34811.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 65:20:@34811.4]
  wire  regs_109_io_enable; // @[RegFile.scala 65:20:@34811.4]
  wire  regs_110_clock; // @[RegFile.scala 65:20:@34825.4]
  wire  regs_110_reset; // @[RegFile.scala 65:20:@34825.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 65:20:@34825.4]
  wire  regs_110_io_reset; // @[RegFile.scala 65:20:@34825.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 65:20:@34825.4]
  wire  regs_110_io_enable; // @[RegFile.scala 65:20:@34825.4]
  wire  regs_111_clock; // @[RegFile.scala 65:20:@34839.4]
  wire  regs_111_reset; // @[RegFile.scala 65:20:@34839.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 65:20:@34839.4]
  wire  regs_111_io_reset; // @[RegFile.scala 65:20:@34839.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 65:20:@34839.4]
  wire  regs_111_io_enable; // @[RegFile.scala 65:20:@34839.4]
  wire  regs_112_clock; // @[RegFile.scala 65:20:@34853.4]
  wire  regs_112_reset; // @[RegFile.scala 65:20:@34853.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 65:20:@34853.4]
  wire  regs_112_io_reset; // @[RegFile.scala 65:20:@34853.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 65:20:@34853.4]
  wire  regs_112_io_enable; // @[RegFile.scala 65:20:@34853.4]
  wire  regs_113_clock; // @[RegFile.scala 65:20:@34867.4]
  wire  regs_113_reset; // @[RegFile.scala 65:20:@34867.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 65:20:@34867.4]
  wire  regs_113_io_reset; // @[RegFile.scala 65:20:@34867.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 65:20:@34867.4]
  wire  regs_113_io_enable; // @[RegFile.scala 65:20:@34867.4]
  wire  regs_114_clock; // @[RegFile.scala 65:20:@34881.4]
  wire  regs_114_reset; // @[RegFile.scala 65:20:@34881.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 65:20:@34881.4]
  wire  regs_114_io_reset; // @[RegFile.scala 65:20:@34881.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 65:20:@34881.4]
  wire  regs_114_io_enable; // @[RegFile.scala 65:20:@34881.4]
  wire  regs_115_clock; // @[RegFile.scala 65:20:@34895.4]
  wire  regs_115_reset; // @[RegFile.scala 65:20:@34895.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 65:20:@34895.4]
  wire  regs_115_io_reset; // @[RegFile.scala 65:20:@34895.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 65:20:@34895.4]
  wire  regs_115_io_enable; // @[RegFile.scala 65:20:@34895.4]
  wire  regs_116_clock; // @[RegFile.scala 65:20:@34909.4]
  wire  regs_116_reset; // @[RegFile.scala 65:20:@34909.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 65:20:@34909.4]
  wire  regs_116_io_reset; // @[RegFile.scala 65:20:@34909.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 65:20:@34909.4]
  wire  regs_116_io_enable; // @[RegFile.scala 65:20:@34909.4]
  wire  regs_117_clock; // @[RegFile.scala 65:20:@34923.4]
  wire  regs_117_reset; // @[RegFile.scala 65:20:@34923.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 65:20:@34923.4]
  wire  regs_117_io_reset; // @[RegFile.scala 65:20:@34923.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 65:20:@34923.4]
  wire  regs_117_io_enable; // @[RegFile.scala 65:20:@34923.4]
  wire  regs_118_clock; // @[RegFile.scala 65:20:@34937.4]
  wire  regs_118_reset; // @[RegFile.scala 65:20:@34937.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 65:20:@34937.4]
  wire  regs_118_io_reset; // @[RegFile.scala 65:20:@34937.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 65:20:@34937.4]
  wire  regs_118_io_enable; // @[RegFile.scala 65:20:@34937.4]
  wire  regs_119_clock; // @[RegFile.scala 65:20:@34951.4]
  wire  regs_119_reset; // @[RegFile.scala 65:20:@34951.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 65:20:@34951.4]
  wire  regs_119_io_reset; // @[RegFile.scala 65:20:@34951.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 65:20:@34951.4]
  wire  regs_119_io_enable; // @[RegFile.scala 65:20:@34951.4]
  wire  regs_120_clock; // @[RegFile.scala 65:20:@34965.4]
  wire  regs_120_reset; // @[RegFile.scala 65:20:@34965.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 65:20:@34965.4]
  wire  regs_120_io_reset; // @[RegFile.scala 65:20:@34965.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 65:20:@34965.4]
  wire  regs_120_io_enable; // @[RegFile.scala 65:20:@34965.4]
  wire  regs_121_clock; // @[RegFile.scala 65:20:@34979.4]
  wire  regs_121_reset; // @[RegFile.scala 65:20:@34979.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 65:20:@34979.4]
  wire  regs_121_io_reset; // @[RegFile.scala 65:20:@34979.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 65:20:@34979.4]
  wire  regs_121_io_enable; // @[RegFile.scala 65:20:@34979.4]
  wire  regs_122_clock; // @[RegFile.scala 65:20:@34993.4]
  wire  regs_122_reset; // @[RegFile.scala 65:20:@34993.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 65:20:@34993.4]
  wire  regs_122_io_reset; // @[RegFile.scala 65:20:@34993.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 65:20:@34993.4]
  wire  regs_122_io_enable; // @[RegFile.scala 65:20:@34993.4]
  wire  regs_123_clock; // @[RegFile.scala 65:20:@35007.4]
  wire  regs_123_reset; // @[RegFile.scala 65:20:@35007.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 65:20:@35007.4]
  wire  regs_123_io_reset; // @[RegFile.scala 65:20:@35007.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 65:20:@35007.4]
  wire  regs_123_io_enable; // @[RegFile.scala 65:20:@35007.4]
  wire  regs_124_clock; // @[RegFile.scala 65:20:@35021.4]
  wire  regs_124_reset; // @[RegFile.scala 65:20:@35021.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 65:20:@35021.4]
  wire  regs_124_io_reset; // @[RegFile.scala 65:20:@35021.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 65:20:@35021.4]
  wire  regs_124_io_enable; // @[RegFile.scala 65:20:@35021.4]
  wire  regs_125_clock; // @[RegFile.scala 65:20:@35035.4]
  wire  regs_125_reset; // @[RegFile.scala 65:20:@35035.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 65:20:@35035.4]
  wire  regs_125_io_reset; // @[RegFile.scala 65:20:@35035.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 65:20:@35035.4]
  wire  regs_125_io_enable; // @[RegFile.scala 65:20:@35035.4]
  wire  regs_126_clock; // @[RegFile.scala 65:20:@35049.4]
  wire  regs_126_reset; // @[RegFile.scala 65:20:@35049.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 65:20:@35049.4]
  wire  regs_126_io_reset; // @[RegFile.scala 65:20:@35049.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 65:20:@35049.4]
  wire  regs_126_io_enable; // @[RegFile.scala 65:20:@35049.4]
  wire  regs_127_clock; // @[RegFile.scala 65:20:@35063.4]
  wire  regs_127_reset; // @[RegFile.scala 65:20:@35063.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 65:20:@35063.4]
  wire  regs_127_io_reset; // @[RegFile.scala 65:20:@35063.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 65:20:@35063.4]
  wire  regs_127_io_enable; // @[RegFile.scala 65:20:@35063.4]
  wire  regs_128_clock; // @[RegFile.scala 65:20:@35077.4]
  wire  regs_128_reset; // @[RegFile.scala 65:20:@35077.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 65:20:@35077.4]
  wire  regs_128_io_reset; // @[RegFile.scala 65:20:@35077.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 65:20:@35077.4]
  wire  regs_128_io_enable; // @[RegFile.scala 65:20:@35077.4]
  wire  regs_129_clock; // @[RegFile.scala 65:20:@35091.4]
  wire  regs_129_reset; // @[RegFile.scala 65:20:@35091.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 65:20:@35091.4]
  wire  regs_129_io_reset; // @[RegFile.scala 65:20:@35091.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 65:20:@35091.4]
  wire  regs_129_io_enable; // @[RegFile.scala 65:20:@35091.4]
  wire  regs_130_clock; // @[RegFile.scala 65:20:@35105.4]
  wire  regs_130_reset; // @[RegFile.scala 65:20:@35105.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 65:20:@35105.4]
  wire  regs_130_io_reset; // @[RegFile.scala 65:20:@35105.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 65:20:@35105.4]
  wire  regs_130_io_enable; // @[RegFile.scala 65:20:@35105.4]
  wire  regs_131_clock; // @[RegFile.scala 65:20:@35119.4]
  wire  regs_131_reset; // @[RegFile.scala 65:20:@35119.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 65:20:@35119.4]
  wire  regs_131_io_reset; // @[RegFile.scala 65:20:@35119.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 65:20:@35119.4]
  wire  regs_131_io_enable; // @[RegFile.scala 65:20:@35119.4]
  wire  regs_132_clock; // @[RegFile.scala 65:20:@35133.4]
  wire  regs_132_reset; // @[RegFile.scala 65:20:@35133.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 65:20:@35133.4]
  wire  regs_132_io_reset; // @[RegFile.scala 65:20:@35133.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 65:20:@35133.4]
  wire  regs_132_io_enable; // @[RegFile.scala 65:20:@35133.4]
  wire  regs_133_clock; // @[RegFile.scala 65:20:@35147.4]
  wire  regs_133_reset; // @[RegFile.scala 65:20:@35147.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 65:20:@35147.4]
  wire  regs_133_io_reset; // @[RegFile.scala 65:20:@35147.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 65:20:@35147.4]
  wire  regs_133_io_enable; // @[RegFile.scala 65:20:@35147.4]
  wire  regs_134_clock; // @[RegFile.scala 65:20:@35161.4]
  wire  regs_134_reset; // @[RegFile.scala 65:20:@35161.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 65:20:@35161.4]
  wire  regs_134_io_reset; // @[RegFile.scala 65:20:@35161.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 65:20:@35161.4]
  wire  regs_134_io_enable; // @[RegFile.scala 65:20:@35161.4]
  wire  regs_135_clock; // @[RegFile.scala 65:20:@35175.4]
  wire  regs_135_reset; // @[RegFile.scala 65:20:@35175.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 65:20:@35175.4]
  wire  regs_135_io_reset; // @[RegFile.scala 65:20:@35175.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 65:20:@35175.4]
  wire  regs_135_io_enable; // @[RegFile.scala 65:20:@35175.4]
  wire  regs_136_clock; // @[RegFile.scala 65:20:@35189.4]
  wire  regs_136_reset; // @[RegFile.scala 65:20:@35189.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 65:20:@35189.4]
  wire  regs_136_io_reset; // @[RegFile.scala 65:20:@35189.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 65:20:@35189.4]
  wire  regs_136_io_enable; // @[RegFile.scala 65:20:@35189.4]
  wire  regs_137_clock; // @[RegFile.scala 65:20:@35203.4]
  wire  regs_137_reset; // @[RegFile.scala 65:20:@35203.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 65:20:@35203.4]
  wire  regs_137_io_reset; // @[RegFile.scala 65:20:@35203.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 65:20:@35203.4]
  wire  regs_137_io_enable; // @[RegFile.scala 65:20:@35203.4]
  wire  regs_138_clock; // @[RegFile.scala 65:20:@35217.4]
  wire  regs_138_reset; // @[RegFile.scala 65:20:@35217.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 65:20:@35217.4]
  wire  regs_138_io_reset; // @[RegFile.scala 65:20:@35217.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 65:20:@35217.4]
  wire  regs_138_io_enable; // @[RegFile.scala 65:20:@35217.4]
  wire  regs_139_clock; // @[RegFile.scala 65:20:@35231.4]
  wire  regs_139_reset; // @[RegFile.scala 65:20:@35231.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 65:20:@35231.4]
  wire  regs_139_io_reset; // @[RegFile.scala 65:20:@35231.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 65:20:@35231.4]
  wire  regs_139_io_enable; // @[RegFile.scala 65:20:@35231.4]
  wire  regs_140_clock; // @[RegFile.scala 65:20:@35245.4]
  wire  regs_140_reset; // @[RegFile.scala 65:20:@35245.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 65:20:@35245.4]
  wire  regs_140_io_reset; // @[RegFile.scala 65:20:@35245.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 65:20:@35245.4]
  wire  regs_140_io_enable; // @[RegFile.scala 65:20:@35245.4]
  wire  regs_141_clock; // @[RegFile.scala 65:20:@35259.4]
  wire  regs_141_reset; // @[RegFile.scala 65:20:@35259.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 65:20:@35259.4]
  wire  regs_141_io_reset; // @[RegFile.scala 65:20:@35259.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 65:20:@35259.4]
  wire  regs_141_io_enable; // @[RegFile.scala 65:20:@35259.4]
  wire  regs_142_clock; // @[RegFile.scala 65:20:@35273.4]
  wire  regs_142_reset; // @[RegFile.scala 65:20:@35273.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 65:20:@35273.4]
  wire  regs_142_io_reset; // @[RegFile.scala 65:20:@35273.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 65:20:@35273.4]
  wire  regs_142_io_enable; // @[RegFile.scala 65:20:@35273.4]
  wire  regs_143_clock; // @[RegFile.scala 65:20:@35287.4]
  wire  regs_143_reset; // @[RegFile.scala 65:20:@35287.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 65:20:@35287.4]
  wire  regs_143_io_reset; // @[RegFile.scala 65:20:@35287.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 65:20:@35287.4]
  wire  regs_143_io_enable; // @[RegFile.scala 65:20:@35287.4]
  wire  regs_144_clock; // @[RegFile.scala 65:20:@35301.4]
  wire  regs_144_reset; // @[RegFile.scala 65:20:@35301.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 65:20:@35301.4]
  wire  regs_144_io_reset; // @[RegFile.scala 65:20:@35301.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 65:20:@35301.4]
  wire  regs_144_io_enable; // @[RegFile.scala 65:20:@35301.4]
  wire  regs_145_clock; // @[RegFile.scala 65:20:@35315.4]
  wire  regs_145_reset; // @[RegFile.scala 65:20:@35315.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 65:20:@35315.4]
  wire  regs_145_io_reset; // @[RegFile.scala 65:20:@35315.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 65:20:@35315.4]
  wire  regs_145_io_enable; // @[RegFile.scala 65:20:@35315.4]
  wire  regs_146_clock; // @[RegFile.scala 65:20:@35329.4]
  wire  regs_146_reset; // @[RegFile.scala 65:20:@35329.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 65:20:@35329.4]
  wire  regs_146_io_reset; // @[RegFile.scala 65:20:@35329.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 65:20:@35329.4]
  wire  regs_146_io_enable; // @[RegFile.scala 65:20:@35329.4]
  wire  regs_147_clock; // @[RegFile.scala 65:20:@35343.4]
  wire  regs_147_reset; // @[RegFile.scala 65:20:@35343.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 65:20:@35343.4]
  wire  regs_147_io_reset; // @[RegFile.scala 65:20:@35343.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 65:20:@35343.4]
  wire  regs_147_io_enable; // @[RegFile.scala 65:20:@35343.4]
  wire  regs_148_clock; // @[RegFile.scala 65:20:@35357.4]
  wire  regs_148_reset; // @[RegFile.scala 65:20:@35357.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 65:20:@35357.4]
  wire  regs_148_io_reset; // @[RegFile.scala 65:20:@35357.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 65:20:@35357.4]
  wire  regs_148_io_enable; // @[RegFile.scala 65:20:@35357.4]
  wire  regs_149_clock; // @[RegFile.scala 65:20:@35371.4]
  wire  regs_149_reset; // @[RegFile.scala 65:20:@35371.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 65:20:@35371.4]
  wire  regs_149_io_reset; // @[RegFile.scala 65:20:@35371.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 65:20:@35371.4]
  wire  regs_149_io_enable; // @[RegFile.scala 65:20:@35371.4]
  wire  regs_150_clock; // @[RegFile.scala 65:20:@35385.4]
  wire  regs_150_reset; // @[RegFile.scala 65:20:@35385.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 65:20:@35385.4]
  wire  regs_150_io_reset; // @[RegFile.scala 65:20:@35385.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 65:20:@35385.4]
  wire  regs_150_io_enable; // @[RegFile.scala 65:20:@35385.4]
  wire  regs_151_clock; // @[RegFile.scala 65:20:@35399.4]
  wire  regs_151_reset; // @[RegFile.scala 65:20:@35399.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 65:20:@35399.4]
  wire  regs_151_io_reset; // @[RegFile.scala 65:20:@35399.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 65:20:@35399.4]
  wire  regs_151_io_enable; // @[RegFile.scala 65:20:@35399.4]
  wire  regs_152_clock; // @[RegFile.scala 65:20:@35413.4]
  wire  regs_152_reset; // @[RegFile.scala 65:20:@35413.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 65:20:@35413.4]
  wire  regs_152_io_reset; // @[RegFile.scala 65:20:@35413.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 65:20:@35413.4]
  wire  regs_152_io_enable; // @[RegFile.scala 65:20:@35413.4]
  wire  regs_153_clock; // @[RegFile.scala 65:20:@35427.4]
  wire  regs_153_reset; // @[RegFile.scala 65:20:@35427.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 65:20:@35427.4]
  wire  regs_153_io_reset; // @[RegFile.scala 65:20:@35427.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 65:20:@35427.4]
  wire  regs_153_io_enable; // @[RegFile.scala 65:20:@35427.4]
  wire  regs_154_clock; // @[RegFile.scala 65:20:@35441.4]
  wire  regs_154_reset; // @[RegFile.scala 65:20:@35441.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 65:20:@35441.4]
  wire  regs_154_io_reset; // @[RegFile.scala 65:20:@35441.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 65:20:@35441.4]
  wire  regs_154_io_enable; // @[RegFile.scala 65:20:@35441.4]
  wire  regs_155_clock; // @[RegFile.scala 65:20:@35455.4]
  wire  regs_155_reset; // @[RegFile.scala 65:20:@35455.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 65:20:@35455.4]
  wire  regs_155_io_reset; // @[RegFile.scala 65:20:@35455.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 65:20:@35455.4]
  wire  regs_155_io_enable; // @[RegFile.scala 65:20:@35455.4]
  wire  regs_156_clock; // @[RegFile.scala 65:20:@35469.4]
  wire  regs_156_reset; // @[RegFile.scala 65:20:@35469.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 65:20:@35469.4]
  wire  regs_156_io_reset; // @[RegFile.scala 65:20:@35469.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 65:20:@35469.4]
  wire  regs_156_io_enable; // @[RegFile.scala 65:20:@35469.4]
  wire  regs_157_clock; // @[RegFile.scala 65:20:@35483.4]
  wire  regs_157_reset; // @[RegFile.scala 65:20:@35483.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 65:20:@35483.4]
  wire  regs_157_io_reset; // @[RegFile.scala 65:20:@35483.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 65:20:@35483.4]
  wire  regs_157_io_enable; // @[RegFile.scala 65:20:@35483.4]
  wire  regs_158_clock; // @[RegFile.scala 65:20:@35497.4]
  wire  regs_158_reset; // @[RegFile.scala 65:20:@35497.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 65:20:@35497.4]
  wire  regs_158_io_reset; // @[RegFile.scala 65:20:@35497.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 65:20:@35497.4]
  wire  regs_158_io_enable; // @[RegFile.scala 65:20:@35497.4]
  wire  regs_159_clock; // @[RegFile.scala 65:20:@35511.4]
  wire  regs_159_reset; // @[RegFile.scala 65:20:@35511.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 65:20:@35511.4]
  wire  regs_159_io_reset; // @[RegFile.scala 65:20:@35511.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 65:20:@35511.4]
  wire  regs_159_io_enable; // @[RegFile.scala 65:20:@35511.4]
  wire  regs_160_clock; // @[RegFile.scala 65:20:@35525.4]
  wire  regs_160_reset; // @[RegFile.scala 65:20:@35525.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 65:20:@35525.4]
  wire  regs_160_io_reset; // @[RegFile.scala 65:20:@35525.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 65:20:@35525.4]
  wire  regs_160_io_enable; // @[RegFile.scala 65:20:@35525.4]
  wire  regs_161_clock; // @[RegFile.scala 65:20:@35539.4]
  wire  regs_161_reset; // @[RegFile.scala 65:20:@35539.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 65:20:@35539.4]
  wire  regs_161_io_reset; // @[RegFile.scala 65:20:@35539.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 65:20:@35539.4]
  wire  regs_161_io_enable; // @[RegFile.scala 65:20:@35539.4]
  wire  regs_162_clock; // @[RegFile.scala 65:20:@35553.4]
  wire  regs_162_reset; // @[RegFile.scala 65:20:@35553.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 65:20:@35553.4]
  wire  regs_162_io_reset; // @[RegFile.scala 65:20:@35553.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 65:20:@35553.4]
  wire  regs_162_io_enable; // @[RegFile.scala 65:20:@35553.4]
  wire  regs_163_clock; // @[RegFile.scala 65:20:@35567.4]
  wire  regs_163_reset; // @[RegFile.scala 65:20:@35567.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 65:20:@35567.4]
  wire  regs_163_io_reset; // @[RegFile.scala 65:20:@35567.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 65:20:@35567.4]
  wire  regs_163_io_enable; // @[RegFile.scala 65:20:@35567.4]
  wire  regs_164_clock; // @[RegFile.scala 65:20:@35581.4]
  wire  regs_164_reset; // @[RegFile.scala 65:20:@35581.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 65:20:@35581.4]
  wire  regs_164_io_reset; // @[RegFile.scala 65:20:@35581.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 65:20:@35581.4]
  wire  regs_164_io_enable; // @[RegFile.scala 65:20:@35581.4]
  wire  regs_165_clock; // @[RegFile.scala 65:20:@35595.4]
  wire  regs_165_reset; // @[RegFile.scala 65:20:@35595.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 65:20:@35595.4]
  wire  regs_165_io_reset; // @[RegFile.scala 65:20:@35595.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 65:20:@35595.4]
  wire  regs_165_io_enable; // @[RegFile.scala 65:20:@35595.4]
  wire  regs_166_clock; // @[RegFile.scala 65:20:@35609.4]
  wire  regs_166_reset; // @[RegFile.scala 65:20:@35609.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 65:20:@35609.4]
  wire  regs_166_io_reset; // @[RegFile.scala 65:20:@35609.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 65:20:@35609.4]
  wire  regs_166_io_enable; // @[RegFile.scala 65:20:@35609.4]
  wire  regs_167_clock; // @[RegFile.scala 65:20:@35623.4]
  wire  regs_167_reset; // @[RegFile.scala 65:20:@35623.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 65:20:@35623.4]
  wire  regs_167_io_reset; // @[RegFile.scala 65:20:@35623.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 65:20:@35623.4]
  wire  regs_167_io_enable; // @[RegFile.scala 65:20:@35623.4]
  wire  regs_168_clock; // @[RegFile.scala 65:20:@35637.4]
  wire  regs_168_reset; // @[RegFile.scala 65:20:@35637.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 65:20:@35637.4]
  wire  regs_168_io_reset; // @[RegFile.scala 65:20:@35637.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 65:20:@35637.4]
  wire  regs_168_io_enable; // @[RegFile.scala 65:20:@35637.4]
  wire  regs_169_clock; // @[RegFile.scala 65:20:@35651.4]
  wire  regs_169_reset; // @[RegFile.scala 65:20:@35651.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 65:20:@35651.4]
  wire  regs_169_io_reset; // @[RegFile.scala 65:20:@35651.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 65:20:@35651.4]
  wire  regs_169_io_enable; // @[RegFile.scala 65:20:@35651.4]
  wire  regs_170_clock; // @[RegFile.scala 65:20:@35665.4]
  wire  regs_170_reset; // @[RegFile.scala 65:20:@35665.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 65:20:@35665.4]
  wire  regs_170_io_reset; // @[RegFile.scala 65:20:@35665.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 65:20:@35665.4]
  wire  regs_170_io_enable; // @[RegFile.scala 65:20:@35665.4]
  wire  regs_171_clock; // @[RegFile.scala 65:20:@35679.4]
  wire  regs_171_reset; // @[RegFile.scala 65:20:@35679.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 65:20:@35679.4]
  wire  regs_171_io_reset; // @[RegFile.scala 65:20:@35679.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 65:20:@35679.4]
  wire  regs_171_io_enable; // @[RegFile.scala 65:20:@35679.4]
  wire  regs_172_clock; // @[RegFile.scala 65:20:@35693.4]
  wire  regs_172_reset; // @[RegFile.scala 65:20:@35693.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 65:20:@35693.4]
  wire  regs_172_io_reset; // @[RegFile.scala 65:20:@35693.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 65:20:@35693.4]
  wire  regs_172_io_enable; // @[RegFile.scala 65:20:@35693.4]
  wire  regs_173_clock; // @[RegFile.scala 65:20:@35707.4]
  wire  regs_173_reset; // @[RegFile.scala 65:20:@35707.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 65:20:@35707.4]
  wire  regs_173_io_reset; // @[RegFile.scala 65:20:@35707.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 65:20:@35707.4]
  wire  regs_173_io_enable; // @[RegFile.scala 65:20:@35707.4]
  wire  regs_174_clock; // @[RegFile.scala 65:20:@35721.4]
  wire  regs_174_reset; // @[RegFile.scala 65:20:@35721.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 65:20:@35721.4]
  wire  regs_174_io_reset; // @[RegFile.scala 65:20:@35721.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 65:20:@35721.4]
  wire  regs_174_io_enable; // @[RegFile.scala 65:20:@35721.4]
  wire  regs_175_clock; // @[RegFile.scala 65:20:@35735.4]
  wire  regs_175_reset; // @[RegFile.scala 65:20:@35735.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 65:20:@35735.4]
  wire  regs_175_io_reset; // @[RegFile.scala 65:20:@35735.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 65:20:@35735.4]
  wire  regs_175_io_enable; // @[RegFile.scala 65:20:@35735.4]
  wire  regs_176_clock; // @[RegFile.scala 65:20:@35749.4]
  wire  regs_176_reset; // @[RegFile.scala 65:20:@35749.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 65:20:@35749.4]
  wire  regs_176_io_reset; // @[RegFile.scala 65:20:@35749.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 65:20:@35749.4]
  wire  regs_176_io_enable; // @[RegFile.scala 65:20:@35749.4]
  wire  regs_177_clock; // @[RegFile.scala 65:20:@35763.4]
  wire  regs_177_reset; // @[RegFile.scala 65:20:@35763.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 65:20:@35763.4]
  wire  regs_177_io_reset; // @[RegFile.scala 65:20:@35763.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 65:20:@35763.4]
  wire  regs_177_io_enable; // @[RegFile.scala 65:20:@35763.4]
  wire  regs_178_clock; // @[RegFile.scala 65:20:@35777.4]
  wire  regs_178_reset; // @[RegFile.scala 65:20:@35777.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 65:20:@35777.4]
  wire  regs_178_io_reset; // @[RegFile.scala 65:20:@35777.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 65:20:@35777.4]
  wire  regs_178_io_enable; // @[RegFile.scala 65:20:@35777.4]
  wire  regs_179_clock; // @[RegFile.scala 65:20:@35791.4]
  wire  regs_179_reset; // @[RegFile.scala 65:20:@35791.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 65:20:@35791.4]
  wire  regs_179_io_reset; // @[RegFile.scala 65:20:@35791.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 65:20:@35791.4]
  wire  regs_179_io_enable; // @[RegFile.scala 65:20:@35791.4]
  wire  regs_180_clock; // @[RegFile.scala 65:20:@35805.4]
  wire  regs_180_reset; // @[RegFile.scala 65:20:@35805.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 65:20:@35805.4]
  wire  regs_180_io_reset; // @[RegFile.scala 65:20:@35805.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 65:20:@35805.4]
  wire  regs_180_io_enable; // @[RegFile.scala 65:20:@35805.4]
  wire  regs_181_clock; // @[RegFile.scala 65:20:@35819.4]
  wire  regs_181_reset; // @[RegFile.scala 65:20:@35819.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 65:20:@35819.4]
  wire  regs_181_io_reset; // @[RegFile.scala 65:20:@35819.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 65:20:@35819.4]
  wire  regs_181_io_enable; // @[RegFile.scala 65:20:@35819.4]
  wire  regs_182_clock; // @[RegFile.scala 65:20:@35833.4]
  wire  regs_182_reset; // @[RegFile.scala 65:20:@35833.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 65:20:@35833.4]
  wire  regs_182_io_reset; // @[RegFile.scala 65:20:@35833.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 65:20:@35833.4]
  wire  regs_182_io_enable; // @[RegFile.scala 65:20:@35833.4]
  wire  regs_183_clock; // @[RegFile.scala 65:20:@35847.4]
  wire  regs_183_reset; // @[RegFile.scala 65:20:@35847.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 65:20:@35847.4]
  wire  regs_183_io_reset; // @[RegFile.scala 65:20:@35847.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 65:20:@35847.4]
  wire  regs_183_io_enable; // @[RegFile.scala 65:20:@35847.4]
  wire  regs_184_clock; // @[RegFile.scala 65:20:@35861.4]
  wire  regs_184_reset; // @[RegFile.scala 65:20:@35861.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 65:20:@35861.4]
  wire  regs_184_io_reset; // @[RegFile.scala 65:20:@35861.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 65:20:@35861.4]
  wire  regs_184_io_enable; // @[RegFile.scala 65:20:@35861.4]
  wire  regs_185_clock; // @[RegFile.scala 65:20:@35875.4]
  wire  regs_185_reset; // @[RegFile.scala 65:20:@35875.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 65:20:@35875.4]
  wire  regs_185_io_reset; // @[RegFile.scala 65:20:@35875.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 65:20:@35875.4]
  wire  regs_185_io_enable; // @[RegFile.scala 65:20:@35875.4]
  wire  regs_186_clock; // @[RegFile.scala 65:20:@35889.4]
  wire  regs_186_reset; // @[RegFile.scala 65:20:@35889.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 65:20:@35889.4]
  wire  regs_186_io_reset; // @[RegFile.scala 65:20:@35889.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 65:20:@35889.4]
  wire  regs_186_io_enable; // @[RegFile.scala 65:20:@35889.4]
  wire  regs_187_clock; // @[RegFile.scala 65:20:@35903.4]
  wire  regs_187_reset; // @[RegFile.scala 65:20:@35903.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 65:20:@35903.4]
  wire  regs_187_io_reset; // @[RegFile.scala 65:20:@35903.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 65:20:@35903.4]
  wire  regs_187_io_enable; // @[RegFile.scala 65:20:@35903.4]
  wire  regs_188_clock; // @[RegFile.scala 65:20:@35917.4]
  wire  regs_188_reset; // @[RegFile.scala 65:20:@35917.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 65:20:@35917.4]
  wire  regs_188_io_reset; // @[RegFile.scala 65:20:@35917.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 65:20:@35917.4]
  wire  regs_188_io_enable; // @[RegFile.scala 65:20:@35917.4]
  wire  regs_189_clock; // @[RegFile.scala 65:20:@35931.4]
  wire  regs_189_reset; // @[RegFile.scala 65:20:@35931.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 65:20:@35931.4]
  wire  regs_189_io_reset; // @[RegFile.scala 65:20:@35931.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 65:20:@35931.4]
  wire  regs_189_io_enable; // @[RegFile.scala 65:20:@35931.4]
  wire  regs_190_clock; // @[RegFile.scala 65:20:@35945.4]
  wire  regs_190_reset; // @[RegFile.scala 65:20:@35945.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 65:20:@35945.4]
  wire  regs_190_io_reset; // @[RegFile.scala 65:20:@35945.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 65:20:@35945.4]
  wire  regs_190_io_enable; // @[RegFile.scala 65:20:@35945.4]
  wire  regs_191_clock; // @[RegFile.scala 65:20:@35959.4]
  wire  regs_191_reset; // @[RegFile.scala 65:20:@35959.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 65:20:@35959.4]
  wire  regs_191_io_reset; // @[RegFile.scala 65:20:@35959.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 65:20:@35959.4]
  wire  regs_191_io_enable; // @[RegFile.scala 65:20:@35959.4]
  wire  regs_192_clock; // @[RegFile.scala 65:20:@35973.4]
  wire  regs_192_reset; // @[RegFile.scala 65:20:@35973.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 65:20:@35973.4]
  wire  regs_192_io_reset; // @[RegFile.scala 65:20:@35973.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 65:20:@35973.4]
  wire  regs_192_io_enable; // @[RegFile.scala 65:20:@35973.4]
  wire  regs_193_clock; // @[RegFile.scala 65:20:@35987.4]
  wire  regs_193_reset; // @[RegFile.scala 65:20:@35987.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 65:20:@35987.4]
  wire  regs_193_io_reset; // @[RegFile.scala 65:20:@35987.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 65:20:@35987.4]
  wire  regs_193_io_enable; // @[RegFile.scala 65:20:@35987.4]
  wire  regs_194_clock; // @[RegFile.scala 65:20:@36001.4]
  wire  regs_194_reset; // @[RegFile.scala 65:20:@36001.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 65:20:@36001.4]
  wire  regs_194_io_reset; // @[RegFile.scala 65:20:@36001.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 65:20:@36001.4]
  wire  regs_194_io_enable; // @[RegFile.scala 65:20:@36001.4]
  wire  regs_195_clock; // @[RegFile.scala 65:20:@36015.4]
  wire  regs_195_reset; // @[RegFile.scala 65:20:@36015.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 65:20:@36015.4]
  wire  regs_195_io_reset; // @[RegFile.scala 65:20:@36015.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 65:20:@36015.4]
  wire  regs_195_io_enable; // @[RegFile.scala 65:20:@36015.4]
  wire  regs_196_clock; // @[RegFile.scala 65:20:@36029.4]
  wire  regs_196_reset; // @[RegFile.scala 65:20:@36029.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 65:20:@36029.4]
  wire  regs_196_io_reset; // @[RegFile.scala 65:20:@36029.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 65:20:@36029.4]
  wire  regs_196_io_enable; // @[RegFile.scala 65:20:@36029.4]
  wire  regs_197_clock; // @[RegFile.scala 65:20:@36043.4]
  wire  regs_197_reset; // @[RegFile.scala 65:20:@36043.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 65:20:@36043.4]
  wire  regs_197_io_reset; // @[RegFile.scala 65:20:@36043.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 65:20:@36043.4]
  wire  regs_197_io_enable; // @[RegFile.scala 65:20:@36043.4]
  wire  regs_198_clock; // @[RegFile.scala 65:20:@36057.4]
  wire  regs_198_reset; // @[RegFile.scala 65:20:@36057.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 65:20:@36057.4]
  wire  regs_198_io_reset; // @[RegFile.scala 65:20:@36057.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 65:20:@36057.4]
  wire  regs_198_io_enable; // @[RegFile.scala 65:20:@36057.4]
  wire  regs_199_clock; // @[RegFile.scala 65:20:@36071.4]
  wire  regs_199_reset; // @[RegFile.scala 65:20:@36071.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 65:20:@36071.4]
  wire  regs_199_io_reset; // @[RegFile.scala 65:20:@36071.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 65:20:@36071.4]
  wire  regs_199_io_enable; // @[RegFile.scala 65:20:@36071.4]
  wire  regs_200_clock; // @[RegFile.scala 65:20:@36085.4]
  wire  regs_200_reset; // @[RegFile.scala 65:20:@36085.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 65:20:@36085.4]
  wire  regs_200_io_reset; // @[RegFile.scala 65:20:@36085.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 65:20:@36085.4]
  wire  regs_200_io_enable; // @[RegFile.scala 65:20:@36085.4]
  wire  regs_201_clock; // @[RegFile.scala 65:20:@36099.4]
  wire  regs_201_reset; // @[RegFile.scala 65:20:@36099.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 65:20:@36099.4]
  wire  regs_201_io_reset; // @[RegFile.scala 65:20:@36099.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 65:20:@36099.4]
  wire  regs_201_io_enable; // @[RegFile.scala 65:20:@36099.4]
  wire  regs_202_clock; // @[RegFile.scala 65:20:@36113.4]
  wire  regs_202_reset; // @[RegFile.scala 65:20:@36113.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 65:20:@36113.4]
  wire  regs_202_io_reset; // @[RegFile.scala 65:20:@36113.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 65:20:@36113.4]
  wire  regs_202_io_enable; // @[RegFile.scala 65:20:@36113.4]
  wire  regs_203_clock; // @[RegFile.scala 65:20:@36127.4]
  wire  regs_203_reset; // @[RegFile.scala 65:20:@36127.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 65:20:@36127.4]
  wire  regs_203_io_reset; // @[RegFile.scala 65:20:@36127.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 65:20:@36127.4]
  wire  regs_203_io_enable; // @[RegFile.scala 65:20:@36127.4]
  wire  regs_204_clock; // @[RegFile.scala 65:20:@36141.4]
  wire  regs_204_reset; // @[RegFile.scala 65:20:@36141.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 65:20:@36141.4]
  wire  regs_204_io_reset; // @[RegFile.scala 65:20:@36141.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 65:20:@36141.4]
  wire  regs_204_io_enable; // @[RegFile.scala 65:20:@36141.4]
  wire  regs_205_clock; // @[RegFile.scala 65:20:@36155.4]
  wire  regs_205_reset; // @[RegFile.scala 65:20:@36155.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 65:20:@36155.4]
  wire  regs_205_io_reset; // @[RegFile.scala 65:20:@36155.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 65:20:@36155.4]
  wire  regs_205_io_enable; // @[RegFile.scala 65:20:@36155.4]
  wire  regs_206_clock; // @[RegFile.scala 65:20:@36169.4]
  wire  regs_206_reset; // @[RegFile.scala 65:20:@36169.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 65:20:@36169.4]
  wire  regs_206_io_reset; // @[RegFile.scala 65:20:@36169.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 65:20:@36169.4]
  wire  regs_206_io_enable; // @[RegFile.scala 65:20:@36169.4]
  wire  regs_207_clock; // @[RegFile.scala 65:20:@36183.4]
  wire  regs_207_reset; // @[RegFile.scala 65:20:@36183.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 65:20:@36183.4]
  wire  regs_207_io_reset; // @[RegFile.scala 65:20:@36183.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 65:20:@36183.4]
  wire  regs_207_io_enable; // @[RegFile.scala 65:20:@36183.4]
  wire  regs_208_clock; // @[RegFile.scala 65:20:@36197.4]
  wire  regs_208_reset; // @[RegFile.scala 65:20:@36197.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 65:20:@36197.4]
  wire  regs_208_io_reset; // @[RegFile.scala 65:20:@36197.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 65:20:@36197.4]
  wire  regs_208_io_enable; // @[RegFile.scala 65:20:@36197.4]
  wire  regs_209_clock; // @[RegFile.scala 65:20:@36211.4]
  wire  regs_209_reset; // @[RegFile.scala 65:20:@36211.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 65:20:@36211.4]
  wire  regs_209_io_reset; // @[RegFile.scala 65:20:@36211.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 65:20:@36211.4]
  wire  regs_209_io_enable; // @[RegFile.scala 65:20:@36211.4]
  wire  regs_210_clock; // @[RegFile.scala 65:20:@36225.4]
  wire  regs_210_reset; // @[RegFile.scala 65:20:@36225.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 65:20:@36225.4]
  wire  regs_210_io_reset; // @[RegFile.scala 65:20:@36225.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 65:20:@36225.4]
  wire  regs_210_io_enable; // @[RegFile.scala 65:20:@36225.4]
  wire  regs_211_clock; // @[RegFile.scala 65:20:@36239.4]
  wire  regs_211_reset; // @[RegFile.scala 65:20:@36239.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 65:20:@36239.4]
  wire  regs_211_io_reset; // @[RegFile.scala 65:20:@36239.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 65:20:@36239.4]
  wire  regs_211_io_enable; // @[RegFile.scala 65:20:@36239.4]
  wire  regs_212_clock; // @[RegFile.scala 65:20:@36253.4]
  wire  regs_212_reset; // @[RegFile.scala 65:20:@36253.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 65:20:@36253.4]
  wire  regs_212_io_reset; // @[RegFile.scala 65:20:@36253.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 65:20:@36253.4]
  wire  regs_212_io_enable; // @[RegFile.scala 65:20:@36253.4]
  wire  regs_213_clock; // @[RegFile.scala 65:20:@36267.4]
  wire  regs_213_reset; // @[RegFile.scala 65:20:@36267.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 65:20:@36267.4]
  wire  regs_213_io_reset; // @[RegFile.scala 65:20:@36267.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 65:20:@36267.4]
  wire  regs_213_io_enable; // @[RegFile.scala 65:20:@36267.4]
  wire  regs_214_clock; // @[RegFile.scala 65:20:@36281.4]
  wire  regs_214_reset; // @[RegFile.scala 65:20:@36281.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 65:20:@36281.4]
  wire  regs_214_io_reset; // @[RegFile.scala 65:20:@36281.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 65:20:@36281.4]
  wire  regs_214_io_enable; // @[RegFile.scala 65:20:@36281.4]
  wire  regs_215_clock; // @[RegFile.scala 65:20:@36295.4]
  wire  regs_215_reset; // @[RegFile.scala 65:20:@36295.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 65:20:@36295.4]
  wire  regs_215_io_reset; // @[RegFile.scala 65:20:@36295.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 65:20:@36295.4]
  wire  regs_215_io_enable; // @[RegFile.scala 65:20:@36295.4]
  wire  regs_216_clock; // @[RegFile.scala 65:20:@36309.4]
  wire  regs_216_reset; // @[RegFile.scala 65:20:@36309.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 65:20:@36309.4]
  wire  regs_216_io_reset; // @[RegFile.scala 65:20:@36309.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 65:20:@36309.4]
  wire  regs_216_io_enable; // @[RegFile.scala 65:20:@36309.4]
  wire  regs_217_clock; // @[RegFile.scala 65:20:@36323.4]
  wire  regs_217_reset; // @[RegFile.scala 65:20:@36323.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 65:20:@36323.4]
  wire  regs_217_io_reset; // @[RegFile.scala 65:20:@36323.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 65:20:@36323.4]
  wire  regs_217_io_enable; // @[RegFile.scala 65:20:@36323.4]
  wire  regs_218_clock; // @[RegFile.scala 65:20:@36337.4]
  wire  regs_218_reset; // @[RegFile.scala 65:20:@36337.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 65:20:@36337.4]
  wire  regs_218_io_reset; // @[RegFile.scala 65:20:@36337.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 65:20:@36337.4]
  wire  regs_218_io_enable; // @[RegFile.scala 65:20:@36337.4]
  wire  regs_219_clock; // @[RegFile.scala 65:20:@36351.4]
  wire  regs_219_reset; // @[RegFile.scala 65:20:@36351.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 65:20:@36351.4]
  wire  regs_219_io_reset; // @[RegFile.scala 65:20:@36351.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 65:20:@36351.4]
  wire  regs_219_io_enable; // @[RegFile.scala 65:20:@36351.4]
  wire  regs_220_clock; // @[RegFile.scala 65:20:@36365.4]
  wire  regs_220_reset; // @[RegFile.scala 65:20:@36365.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 65:20:@36365.4]
  wire  regs_220_io_reset; // @[RegFile.scala 65:20:@36365.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 65:20:@36365.4]
  wire  regs_220_io_enable; // @[RegFile.scala 65:20:@36365.4]
  wire  regs_221_clock; // @[RegFile.scala 65:20:@36379.4]
  wire  regs_221_reset; // @[RegFile.scala 65:20:@36379.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 65:20:@36379.4]
  wire  regs_221_io_reset; // @[RegFile.scala 65:20:@36379.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 65:20:@36379.4]
  wire  regs_221_io_enable; // @[RegFile.scala 65:20:@36379.4]
  wire  regs_222_clock; // @[RegFile.scala 65:20:@36393.4]
  wire  regs_222_reset; // @[RegFile.scala 65:20:@36393.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 65:20:@36393.4]
  wire  regs_222_io_reset; // @[RegFile.scala 65:20:@36393.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 65:20:@36393.4]
  wire  regs_222_io_enable; // @[RegFile.scala 65:20:@36393.4]
  wire  regs_223_clock; // @[RegFile.scala 65:20:@36407.4]
  wire  regs_223_reset; // @[RegFile.scala 65:20:@36407.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 65:20:@36407.4]
  wire  regs_223_io_reset; // @[RegFile.scala 65:20:@36407.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 65:20:@36407.4]
  wire  regs_223_io_enable; // @[RegFile.scala 65:20:@36407.4]
  wire  regs_224_clock; // @[RegFile.scala 65:20:@36421.4]
  wire  regs_224_reset; // @[RegFile.scala 65:20:@36421.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 65:20:@36421.4]
  wire  regs_224_io_reset; // @[RegFile.scala 65:20:@36421.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 65:20:@36421.4]
  wire  regs_224_io_enable; // @[RegFile.scala 65:20:@36421.4]
  wire  regs_225_clock; // @[RegFile.scala 65:20:@36435.4]
  wire  regs_225_reset; // @[RegFile.scala 65:20:@36435.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 65:20:@36435.4]
  wire  regs_225_io_reset; // @[RegFile.scala 65:20:@36435.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 65:20:@36435.4]
  wire  regs_225_io_enable; // @[RegFile.scala 65:20:@36435.4]
  wire  regs_226_clock; // @[RegFile.scala 65:20:@36449.4]
  wire  regs_226_reset; // @[RegFile.scala 65:20:@36449.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 65:20:@36449.4]
  wire  regs_226_io_reset; // @[RegFile.scala 65:20:@36449.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 65:20:@36449.4]
  wire  regs_226_io_enable; // @[RegFile.scala 65:20:@36449.4]
  wire  regs_227_clock; // @[RegFile.scala 65:20:@36463.4]
  wire  regs_227_reset; // @[RegFile.scala 65:20:@36463.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 65:20:@36463.4]
  wire  regs_227_io_reset; // @[RegFile.scala 65:20:@36463.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 65:20:@36463.4]
  wire  regs_227_io_enable; // @[RegFile.scala 65:20:@36463.4]
  wire  regs_228_clock; // @[RegFile.scala 65:20:@36477.4]
  wire  regs_228_reset; // @[RegFile.scala 65:20:@36477.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 65:20:@36477.4]
  wire  regs_228_io_reset; // @[RegFile.scala 65:20:@36477.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 65:20:@36477.4]
  wire  regs_228_io_enable; // @[RegFile.scala 65:20:@36477.4]
  wire  regs_229_clock; // @[RegFile.scala 65:20:@36491.4]
  wire  regs_229_reset; // @[RegFile.scala 65:20:@36491.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 65:20:@36491.4]
  wire  regs_229_io_reset; // @[RegFile.scala 65:20:@36491.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 65:20:@36491.4]
  wire  regs_229_io_enable; // @[RegFile.scala 65:20:@36491.4]
  wire  regs_230_clock; // @[RegFile.scala 65:20:@36505.4]
  wire  regs_230_reset; // @[RegFile.scala 65:20:@36505.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 65:20:@36505.4]
  wire  regs_230_io_reset; // @[RegFile.scala 65:20:@36505.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 65:20:@36505.4]
  wire  regs_230_io_enable; // @[RegFile.scala 65:20:@36505.4]
  wire  regs_231_clock; // @[RegFile.scala 65:20:@36519.4]
  wire  regs_231_reset; // @[RegFile.scala 65:20:@36519.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 65:20:@36519.4]
  wire  regs_231_io_reset; // @[RegFile.scala 65:20:@36519.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 65:20:@36519.4]
  wire  regs_231_io_enable; // @[RegFile.scala 65:20:@36519.4]
  wire  regs_232_clock; // @[RegFile.scala 65:20:@36533.4]
  wire  regs_232_reset; // @[RegFile.scala 65:20:@36533.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 65:20:@36533.4]
  wire  regs_232_io_reset; // @[RegFile.scala 65:20:@36533.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 65:20:@36533.4]
  wire  regs_232_io_enable; // @[RegFile.scala 65:20:@36533.4]
  wire  regs_233_clock; // @[RegFile.scala 65:20:@36547.4]
  wire  regs_233_reset; // @[RegFile.scala 65:20:@36547.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 65:20:@36547.4]
  wire  regs_233_io_reset; // @[RegFile.scala 65:20:@36547.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 65:20:@36547.4]
  wire  regs_233_io_enable; // @[RegFile.scala 65:20:@36547.4]
  wire  regs_234_clock; // @[RegFile.scala 65:20:@36561.4]
  wire  regs_234_reset; // @[RegFile.scala 65:20:@36561.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 65:20:@36561.4]
  wire  regs_234_io_reset; // @[RegFile.scala 65:20:@36561.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 65:20:@36561.4]
  wire  regs_234_io_enable; // @[RegFile.scala 65:20:@36561.4]
  wire  regs_235_clock; // @[RegFile.scala 65:20:@36575.4]
  wire  regs_235_reset; // @[RegFile.scala 65:20:@36575.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 65:20:@36575.4]
  wire  regs_235_io_reset; // @[RegFile.scala 65:20:@36575.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 65:20:@36575.4]
  wire  regs_235_io_enable; // @[RegFile.scala 65:20:@36575.4]
  wire  regs_236_clock; // @[RegFile.scala 65:20:@36589.4]
  wire  regs_236_reset; // @[RegFile.scala 65:20:@36589.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 65:20:@36589.4]
  wire  regs_236_io_reset; // @[RegFile.scala 65:20:@36589.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 65:20:@36589.4]
  wire  regs_236_io_enable; // @[RegFile.scala 65:20:@36589.4]
  wire  regs_237_clock; // @[RegFile.scala 65:20:@36603.4]
  wire  regs_237_reset; // @[RegFile.scala 65:20:@36603.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 65:20:@36603.4]
  wire  regs_237_io_reset; // @[RegFile.scala 65:20:@36603.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 65:20:@36603.4]
  wire  regs_237_io_enable; // @[RegFile.scala 65:20:@36603.4]
  wire  regs_238_clock; // @[RegFile.scala 65:20:@36617.4]
  wire  regs_238_reset; // @[RegFile.scala 65:20:@36617.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 65:20:@36617.4]
  wire  regs_238_io_reset; // @[RegFile.scala 65:20:@36617.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 65:20:@36617.4]
  wire  regs_238_io_enable; // @[RegFile.scala 65:20:@36617.4]
  wire  regs_239_clock; // @[RegFile.scala 65:20:@36631.4]
  wire  regs_239_reset; // @[RegFile.scala 65:20:@36631.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 65:20:@36631.4]
  wire  regs_239_io_reset; // @[RegFile.scala 65:20:@36631.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 65:20:@36631.4]
  wire  regs_239_io_enable; // @[RegFile.scala 65:20:@36631.4]
  wire  regs_240_clock; // @[RegFile.scala 65:20:@36645.4]
  wire  regs_240_reset; // @[RegFile.scala 65:20:@36645.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 65:20:@36645.4]
  wire  regs_240_io_reset; // @[RegFile.scala 65:20:@36645.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 65:20:@36645.4]
  wire  regs_240_io_enable; // @[RegFile.scala 65:20:@36645.4]
  wire  regs_241_clock; // @[RegFile.scala 65:20:@36659.4]
  wire  regs_241_reset; // @[RegFile.scala 65:20:@36659.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 65:20:@36659.4]
  wire  regs_241_io_reset; // @[RegFile.scala 65:20:@36659.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 65:20:@36659.4]
  wire  regs_241_io_enable; // @[RegFile.scala 65:20:@36659.4]
  wire  regs_242_clock; // @[RegFile.scala 65:20:@36673.4]
  wire  regs_242_reset; // @[RegFile.scala 65:20:@36673.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 65:20:@36673.4]
  wire  regs_242_io_reset; // @[RegFile.scala 65:20:@36673.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 65:20:@36673.4]
  wire  regs_242_io_enable; // @[RegFile.scala 65:20:@36673.4]
  wire  regs_243_clock; // @[RegFile.scala 65:20:@36687.4]
  wire  regs_243_reset; // @[RegFile.scala 65:20:@36687.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 65:20:@36687.4]
  wire  regs_243_io_reset; // @[RegFile.scala 65:20:@36687.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 65:20:@36687.4]
  wire  regs_243_io_enable; // @[RegFile.scala 65:20:@36687.4]
  wire  regs_244_clock; // @[RegFile.scala 65:20:@36701.4]
  wire  regs_244_reset; // @[RegFile.scala 65:20:@36701.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 65:20:@36701.4]
  wire  regs_244_io_reset; // @[RegFile.scala 65:20:@36701.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 65:20:@36701.4]
  wire  regs_244_io_enable; // @[RegFile.scala 65:20:@36701.4]
  wire  regs_245_clock; // @[RegFile.scala 65:20:@36715.4]
  wire  regs_245_reset; // @[RegFile.scala 65:20:@36715.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 65:20:@36715.4]
  wire  regs_245_io_reset; // @[RegFile.scala 65:20:@36715.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 65:20:@36715.4]
  wire  regs_245_io_enable; // @[RegFile.scala 65:20:@36715.4]
  wire  regs_246_clock; // @[RegFile.scala 65:20:@36729.4]
  wire  regs_246_reset; // @[RegFile.scala 65:20:@36729.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 65:20:@36729.4]
  wire  regs_246_io_reset; // @[RegFile.scala 65:20:@36729.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 65:20:@36729.4]
  wire  regs_246_io_enable; // @[RegFile.scala 65:20:@36729.4]
  wire  regs_247_clock; // @[RegFile.scala 65:20:@36743.4]
  wire  regs_247_reset; // @[RegFile.scala 65:20:@36743.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 65:20:@36743.4]
  wire  regs_247_io_reset; // @[RegFile.scala 65:20:@36743.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 65:20:@36743.4]
  wire  regs_247_io_enable; // @[RegFile.scala 65:20:@36743.4]
  wire  regs_248_clock; // @[RegFile.scala 65:20:@36757.4]
  wire  regs_248_reset; // @[RegFile.scala 65:20:@36757.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 65:20:@36757.4]
  wire  regs_248_io_reset; // @[RegFile.scala 65:20:@36757.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 65:20:@36757.4]
  wire  regs_248_io_enable; // @[RegFile.scala 65:20:@36757.4]
  wire  regs_249_clock; // @[RegFile.scala 65:20:@36771.4]
  wire  regs_249_reset; // @[RegFile.scala 65:20:@36771.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 65:20:@36771.4]
  wire  regs_249_io_reset; // @[RegFile.scala 65:20:@36771.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 65:20:@36771.4]
  wire  regs_249_io_enable; // @[RegFile.scala 65:20:@36771.4]
  wire  regs_250_clock; // @[RegFile.scala 65:20:@36785.4]
  wire  regs_250_reset; // @[RegFile.scala 65:20:@36785.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 65:20:@36785.4]
  wire  regs_250_io_reset; // @[RegFile.scala 65:20:@36785.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 65:20:@36785.4]
  wire  regs_250_io_enable; // @[RegFile.scala 65:20:@36785.4]
  wire  regs_251_clock; // @[RegFile.scala 65:20:@36799.4]
  wire  regs_251_reset; // @[RegFile.scala 65:20:@36799.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 65:20:@36799.4]
  wire  regs_251_io_reset; // @[RegFile.scala 65:20:@36799.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 65:20:@36799.4]
  wire  regs_251_io_enable; // @[RegFile.scala 65:20:@36799.4]
  wire  regs_252_clock; // @[RegFile.scala 65:20:@36813.4]
  wire  regs_252_reset; // @[RegFile.scala 65:20:@36813.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 65:20:@36813.4]
  wire  regs_252_io_reset; // @[RegFile.scala 65:20:@36813.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 65:20:@36813.4]
  wire  regs_252_io_enable; // @[RegFile.scala 65:20:@36813.4]
  wire  regs_253_clock; // @[RegFile.scala 65:20:@36827.4]
  wire  regs_253_reset; // @[RegFile.scala 65:20:@36827.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 65:20:@36827.4]
  wire  regs_253_io_reset; // @[RegFile.scala 65:20:@36827.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 65:20:@36827.4]
  wire  regs_253_io_enable; // @[RegFile.scala 65:20:@36827.4]
  wire  regs_254_clock; // @[RegFile.scala 65:20:@36841.4]
  wire  regs_254_reset; // @[RegFile.scala 65:20:@36841.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 65:20:@36841.4]
  wire  regs_254_io_reset; // @[RegFile.scala 65:20:@36841.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 65:20:@36841.4]
  wire  regs_254_io_enable; // @[RegFile.scala 65:20:@36841.4]
  wire  regs_255_clock; // @[RegFile.scala 65:20:@36855.4]
  wire  regs_255_reset; // @[RegFile.scala 65:20:@36855.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 65:20:@36855.4]
  wire  regs_255_io_reset; // @[RegFile.scala 65:20:@36855.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 65:20:@36855.4]
  wire  regs_255_io_enable; // @[RegFile.scala 65:20:@36855.4]
  wire  regs_256_clock; // @[RegFile.scala 65:20:@36869.4]
  wire  regs_256_reset; // @[RegFile.scala 65:20:@36869.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 65:20:@36869.4]
  wire  regs_256_io_reset; // @[RegFile.scala 65:20:@36869.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 65:20:@36869.4]
  wire  regs_256_io_enable; // @[RegFile.scala 65:20:@36869.4]
  wire  regs_257_clock; // @[RegFile.scala 65:20:@36883.4]
  wire  regs_257_reset; // @[RegFile.scala 65:20:@36883.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 65:20:@36883.4]
  wire  regs_257_io_reset; // @[RegFile.scala 65:20:@36883.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 65:20:@36883.4]
  wire  regs_257_io_enable; // @[RegFile.scala 65:20:@36883.4]
  wire  regs_258_clock; // @[RegFile.scala 65:20:@36897.4]
  wire  regs_258_reset; // @[RegFile.scala 65:20:@36897.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 65:20:@36897.4]
  wire  regs_258_io_reset; // @[RegFile.scala 65:20:@36897.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 65:20:@36897.4]
  wire  regs_258_io_enable; // @[RegFile.scala 65:20:@36897.4]
  wire  regs_259_clock; // @[RegFile.scala 65:20:@36911.4]
  wire  regs_259_reset; // @[RegFile.scala 65:20:@36911.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 65:20:@36911.4]
  wire  regs_259_io_reset; // @[RegFile.scala 65:20:@36911.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 65:20:@36911.4]
  wire  regs_259_io_enable; // @[RegFile.scala 65:20:@36911.4]
  wire  regs_260_clock; // @[RegFile.scala 65:20:@36925.4]
  wire  regs_260_reset; // @[RegFile.scala 65:20:@36925.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 65:20:@36925.4]
  wire  regs_260_io_reset; // @[RegFile.scala 65:20:@36925.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 65:20:@36925.4]
  wire  regs_260_io_enable; // @[RegFile.scala 65:20:@36925.4]
  wire  regs_261_clock; // @[RegFile.scala 65:20:@36939.4]
  wire  regs_261_reset; // @[RegFile.scala 65:20:@36939.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 65:20:@36939.4]
  wire  regs_261_io_reset; // @[RegFile.scala 65:20:@36939.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 65:20:@36939.4]
  wire  regs_261_io_enable; // @[RegFile.scala 65:20:@36939.4]
  wire  regs_262_clock; // @[RegFile.scala 65:20:@36953.4]
  wire  regs_262_reset; // @[RegFile.scala 65:20:@36953.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 65:20:@36953.4]
  wire  regs_262_io_reset; // @[RegFile.scala 65:20:@36953.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 65:20:@36953.4]
  wire  regs_262_io_enable; // @[RegFile.scala 65:20:@36953.4]
  wire  regs_263_clock; // @[RegFile.scala 65:20:@36967.4]
  wire  regs_263_reset; // @[RegFile.scala 65:20:@36967.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 65:20:@36967.4]
  wire  regs_263_io_reset; // @[RegFile.scala 65:20:@36967.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 65:20:@36967.4]
  wire  regs_263_io_enable; // @[RegFile.scala 65:20:@36967.4]
  wire  regs_264_clock; // @[RegFile.scala 65:20:@36981.4]
  wire  regs_264_reset; // @[RegFile.scala 65:20:@36981.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 65:20:@36981.4]
  wire  regs_264_io_reset; // @[RegFile.scala 65:20:@36981.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 65:20:@36981.4]
  wire  regs_264_io_enable; // @[RegFile.scala 65:20:@36981.4]
  wire  regs_265_clock; // @[RegFile.scala 65:20:@36995.4]
  wire  regs_265_reset; // @[RegFile.scala 65:20:@36995.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 65:20:@36995.4]
  wire  regs_265_io_reset; // @[RegFile.scala 65:20:@36995.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 65:20:@36995.4]
  wire  regs_265_io_enable; // @[RegFile.scala 65:20:@36995.4]
  wire  regs_266_clock; // @[RegFile.scala 65:20:@37009.4]
  wire  regs_266_reset; // @[RegFile.scala 65:20:@37009.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 65:20:@37009.4]
  wire  regs_266_io_reset; // @[RegFile.scala 65:20:@37009.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 65:20:@37009.4]
  wire  regs_266_io_enable; // @[RegFile.scala 65:20:@37009.4]
  wire  regs_267_clock; // @[RegFile.scala 65:20:@37023.4]
  wire  regs_267_reset; // @[RegFile.scala 65:20:@37023.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 65:20:@37023.4]
  wire  regs_267_io_reset; // @[RegFile.scala 65:20:@37023.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 65:20:@37023.4]
  wire  regs_267_io_enable; // @[RegFile.scala 65:20:@37023.4]
  wire  regs_268_clock; // @[RegFile.scala 65:20:@37037.4]
  wire  regs_268_reset; // @[RegFile.scala 65:20:@37037.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 65:20:@37037.4]
  wire  regs_268_io_reset; // @[RegFile.scala 65:20:@37037.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 65:20:@37037.4]
  wire  regs_268_io_enable; // @[RegFile.scala 65:20:@37037.4]
  wire  regs_269_clock; // @[RegFile.scala 65:20:@37051.4]
  wire  regs_269_reset; // @[RegFile.scala 65:20:@37051.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 65:20:@37051.4]
  wire  regs_269_io_reset; // @[RegFile.scala 65:20:@37051.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 65:20:@37051.4]
  wire  regs_269_io_enable; // @[RegFile.scala 65:20:@37051.4]
  wire  regs_270_clock; // @[RegFile.scala 65:20:@37065.4]
  wire  regs_270_reset; // @[RegFile.scala 65:20:@37065.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 65:20:@37065.4]
  wire  regs_270_io_reset; // @[RegFile.scala 65:20:@37065.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 65:20:@37065.4]
  wire  regs_270_io_enable; // @[RegFile.scala 65:20:@37065.4]
  wire  regs_271_clock; // @[RegFile.scala 65:20:@37079.4]
  wire  regs_271_reset; // @[RegFile.scala 65:20:@37079.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 65:20:@37079.4]
  wire  regs_271_io_reset; // @[RegFile.scala 65:20:@37079.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 65:20:@37079.4]
  wire  regs_271_io_enable; // @[RegFile.scala 65:20:@37079.4]
  wire  regs_272_clock; // @[RegFile.scala 65:20:@37093.4]
  wire  regs_272_reset; // @[RegFile.scala 65:20:@37093.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 65:20:@37093.4]
  wire  regs_272_io_reset; // @[RegFile.scala 65:20:@37093.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 65:20:@37093.4]
  wire  regs_272_io_enable; // @[RegFile.scala 65:20:@37093.4]
  wire  regs_273_clock; // @[RegFile.scala 65:20:@37107.4]
  wire  regs_273_reset; // @[RegFile.scala 65:20:@37107.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 65:20:@37107.4]
  wire  regs_273_io_reset; // @[RegFile.scala 65:20:@37107.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 65:20:@37107.4]
  wire  regs_273_io_enable; // @[RegFile.scala 65:20:@37107.4]
  wire  regs_274_clock; // @[RegFile.scala 65:20:@37121.4]
  wire  regs_274_reset; // @[RegFile.scala 65:20:@37121.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 65:20:@37121.4]
  wire  regs_274_io_reset; // @[RegFile.scala 65:20:@37121.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 65:20:@37121.4]
  wire  regs_274_io_enable; // @[RegFile.scala 65:20:@37121.4]
  wire  regs_275_clock; // @[RegFile.scala 65:20:@37135.4]
  wire  regs_275_reset; // @[RegFile.scala 65:20:@37135.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 65:20:@37135.4]
  wire  regs_275_io_reset; // @[RegFile.scala 65:20:@37135.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 65:20:@37135.4]
  wire  regs_275_io_enable; // @[RegFile.scala 65:20:@37135.4]
  wire  regs_276_clock; // @[RegFile.scala 65:20:@37149.4]
  wire  regs_276_reset; // @[RegFile.scala 65:20:@37149.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 65:20:@37149.4]
  wire  regs_276_io_reset; // @[RegFile.scala 65:20:@37149.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 65:20:@37149.4]
  wire  regs_276_io_enable; // @[RegFile.scala 65:20:@37149.4]
  wire  regs_277_clock; // @[RegFile.scala 65:20:@37163.4]
  wire  regs_277_reset; // @[RegFile.scala 65:20:@37163.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 65:20:@37163.4]
  wire  regs_277_io_reset; // @[RegFile.scala 65:20:@37163.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 65:20:@37163.4]
  wire  regs_277_io_enable; // @[RegFile.scala 65:20:@37163.4]
  wire  regs_278_clock; // @[RegFile.scala 65:20:@37177.4]
  wire  regs_278_reset; // @[RegFile.scala 65:20:@37177.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 65:20:@37177.4]
  wire  regs_278_io_reset; // @[RegFile.scala 65:20:@37177.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 65:20:@37177.4]
  wire  regs_278_io_enable; // @[RegFile.scala 65:20:@37177.4]
  wire  regs_279_clock; // @[RegFile.scala 65:20:@37191.4]
  wire  regs_279_reset; // @[RegFile.scala 65:20:@37191.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 65:20:@37191.4]
  wire  regs_279_io_reset; // @[RegFile.scala 65:20:@37191.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 65:20:@37191.4]
  wire  regs_279_io_enable; // @[RegFile.scala 65:20:@37191.4]
  wire  regs_280_clock; // @[RegFile.scala 65:20:@37205.4]
  wire  regs_280_reset; // @[RegFile.scala 65:20:@37205.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 65:20:@37205.4]
  wire  regs_280_io_reset; // @[RegFile.scala 65:20:@37205.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 65:20:@37205.4]
  wire  regs_280_io_enable; // @[RegFile.scala 65:20:@37205.4]
  wire  regs_281_clock; // @[RegFile.scala 65:20:@37219.4]
  wire  regs_281_reset; // @[RegFile.scala 65:20:@37219.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 65:20:@37219.4]
  wire  regs_281_io_reset; // @[RegFile.scala 65:20:@37219.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 65:20:@37219.4]
  wire  regs_281_io_enable; // @[RegFile.scala 65:20:@37219.4]
  wire  regs_282_clock; // @[RegFile.scala 65:20:@37233.4]
  wire  regs_282_reset; // @[RegFile.scala 65:20:@37233.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 65:20:@37233.4]
  wire  regs_282_io_reset; // @[RegFile.scala 65:20:@37233.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 65:20:@37233.4]
  wire  regs_282_io_enable; // @[RegFile.scala 65:20:@37233.4]
  wire  regs_283_clock; // @[RegFile.scala 65:20:@37247.4]
  wire  regs_283_reset; // @[RegFile.scala 65:20:@37247.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 65:20:@37247.4]
  wire  regs_283_io_reset; // @[RegFile.scala 65:20:@37247.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 65:20:@37247.4]
  wire  regs_283_io_enable; // @[RegFile.scala 65:20:@37247.4]
  wire  regs_284_clock; // @[RegFile.scala 65:20:@37261.4]
  wire  regs_284_reset; // @[RegFile.scala 65:20:@37261.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 65:20:@37261.4]
  wire  regs_284_io_reset; // @[RegFile.scala 65:20:@37261.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 65:20:@37261.4]
  wire  regs_284_io_enable; // @[RegFile.scala 65:20:@37261.4]
  wire  regs_285_clock; // @[RegFile.scala 65:20:@37275.4]
  wire  regs_285_reset; // @[RegFile.scala 65:20:@37275.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 65:20:@37275.4]
  wire  regs_285_io_reset; // @[RegFile.scala 65:20:@37275.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 65:20:@37275.4]
  wire  regs_285_io_enable; // @[RegFile.scala 65:20:@37275.4]
  wire  regs_286_clock; // @[RegFile.scala 65:20:@37289.4]
  wire  regs_286_reset; // @[RegFile.scala 65:20:@37289.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 65:20:@37289.4]
  wire  regs_286_io_reset; // @[RegFile.scala 65:20:@37289.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 65:20:@37289.4]
  wire  regs_286_io_enable; // @[RegFile.scala 65:20:@37289.4]
  wire  regs_287_clock; // @[RegFile.scala 65:20:@37303.4]
  wire  regs_287_reset; // @[RegFile.scala 65:20:@37303.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 65:20:@37303.4]
  wire  regs_287_io_reset; // @[RegFile.scala 65:20:@37303.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 65:20:@37303.4]
  wire  regs_287_io_enable; // @[RegFile.scala 65:20:@37303.4]
  wire  regs_288_clock; // @[RegFile.scala 65:20:@37317.4]
  wire  regs_288_reset; // @[RegFile.scala 65:20:@37317.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 65:20:@37317.4]
  wire  regs_288_io_reset; // @[RegFile.scala 65:20:@37317.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 65:20:@37317.4]
  wire  regs_288_io_enable; // @[RegFile.scala 65:20:@37317.4]
  wire  regs_289_clock; // @[RegFile.scala 65:20:@37331.4]
  wire  regs_289_reset; // @[RegFile.scala 65:20:@37331.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 65:20:@37331.4]
  wire  regs_289_io_reset; // @[RegFile.scala 65:20:@37331.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 65:20:@37331.4]
  wire  regs_289_io_enable; // @[RegFile.scala 65:20:@37331.4]
  wire  regs_290_clock; // @[RegFile.scala 65:20:@37345.4]
  wire  regs_290_reset; // @[RegFile.scala 65:20:@37345.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 65:20:@37345.4]
  wire  regs_290_io_reset; // @[RegFile.scala 65:20:@37345.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 65:20:@37345.4]
  wire  regs_290_io_enable; // @[RegFile.scala 65:20:@37345.4]
  wire  regs_291_clock; // @[RegFile.scala 65:20:@37359.4]
  wire  regs_291_reset; // @[RegFile.scala 65:20:@37359.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 65:20:@37359.4]
  wire  regs_291_io_reset; // @[RegFile.scala 65:20:@37359.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 65:20:@37359.4]
  wire  regs_291_io_enable; // @[RegFile.scala 65:20:@37359.4]
  wire  regs_292_clock; // @[RegFile.scala 65:20:@37373.4]
  wire  regs_292_reset; // @[RegFile.scala 65:20:@37373.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 65:20:@37373.4]
  wire  regs_292_io_reset; // @[RegFile.scala 65:20:@37373.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 65:20:@37373.4]
  wire  regs_292_io_enable; // @[RegFile.scala 65:20:@37373.4]
  wire  regs_293_clock; // @[RegFile.scala 65:20:@37387.4]
  wire  regs_293_reset; // @[RegFile.scala 65:20:@37387.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 65:20:@37387.4]
  wire  regs_293_io_reset; // @[RegFile.scala 65:20:@37387.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 65:20:@37387.4]
  wire  regs_293_io_enable; // @[RegFile.scala 65:20:@37387.4]
  wire  regs_294_clock; // @[RegFile.scala 65:20:@37401.4]
  wire  regs_294_reset; // @[RegFile.scala 65:20:@37401.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 65:20:@37401.4]
  wire  regs_294_io_reset; // @[RegFile.scala 65:20:@37401.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 65:20:@37401.4]
  wire  regs_294_io_enable; // @[RegFile.scala 65:20:@37401.4]
  wire  regs_295_clock; // @[RegFile.scala 65:20:@37415.4]
  wire  regs_295_reset; // @[RegFile.scala 65:20:@37415.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 65:20:@37415.4]
  wire  regs_295_io_reset; // @[RegFile.scala 65:20:@37415.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 65:20:@37415.4]
  wire  regs_295_io_enable; // @[RegFile.scala 65:20:@37415.4]
  wire  regs_296_clock; // @[RegFile.scala 65:20:@37429.4]
  wire  regs_296_reset; // @[RegFile.scala 65:20:@37429.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 65:20:@37429.4]
  wire  regs_296_io_reset; // @[RegFile.scala 65:20:@37429.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 65:20:@37429.4]
  wire  regs_296_io_enable; // @[RegFile.scala 65:20:@37429.4]
  wire  regs_297_clock; // @[RegFile.scala 65:20:@37443.4]
  wire  regs_297_reset; // @[RegFile.scala 65:20:@37443.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 65:20:@37443.4]
  wire  regs_297_io_reset; // @[RegFile.scala 65:20:@37443.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 65:20:@37443.4]
  wire  regs_297_io_enable; // @[RegFile.scala 65:20:@37443.4]
  wire  regs_298_clock; // @[RegFile.scala 65:20:@37457.4]
  wire  regs_298_reset; // @[RegFile.scala 65:20:@37457.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 65:20:@37457.4]
  wire  regs_298_io_reset; // @[RegFile.scala 65:20:@37457.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 65:20:@37457.4]
  wire  regs_298_io_enable; // @[RegFile.scala 65:20:@37457.4]
  wire  regs_299_clock; // @[RegFile.scala 65:20:@37471.4]
  wire  regs_299_reset; // @[RegFile.scala 65:20:@37471.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 65:20:@37471.4]
  wire  regs_299_io_reset; // @[RegFile.scala 65:20:@37471.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 65:20:@37471.4]
  wire  regs_299_io_enable; // @[RegFile.scala 65:20:@37471.4]
  wire  regs_300_clock; // @[RegFile.scala 65:20:@37485.4]
  wire  regs_300_reset; // @[RegFile.scala 65:20:@37485.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 65:20:@37485.4]
  wire  regs_300_io_reset; // @[RegFile.scala 65:20:@37485.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 65:20:@37485.4]
  wire  regs_300_io_enable; // @[RegFile.scala 65:20:@37485.4]
  wire  regs_301_clock; // @[RegFile.scala 65:20:@37499.4]
  wire  regs_301_reset; // @[RegFile.scala 65:20:@37499.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 65:20:@37499.4]
  wire  regs_301_io_reset; // @[RegFile.scala 65:20:@37499.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 65:20:@37499.4]
  wire  regs_301_io_enable; // @[RegFile.scala 65:20:@37499.4]
  wire  regs_302_clock; // @[RegFile.scala 65:20:@37513.4]
  wire  regs_302_reset; // @[RegFile.scala 65:20:@37513.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 65:20:@37513.4]
  wire  regs_302_io_reset; // @[RegFile.scala 65:20:@37513.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 65:20:@37513.4]
  wire  regs_302_io_enable; // @[RegFile.scala 65:20:@37513.4]
  wire  regs_303_clock; // @[RegFile.scala 65:20:@37527.4]
  wire  regs_303_reset; // @[RegFile.scala 65:20:@37527.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 65:20:@37527.4]
  wire  regs_303_io_reset; // @[RegFile.scala 65:20:@37527.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 65:20:@37527.4]
  wire  regs_303_io_enable; // @[RegFile.scala 65:20:@37527.4]
  wire  regs_304_clock; // @[RegFile.scala 65:20:@37541.4]
  wire  regs_304_reset; // @[RegFile.scala 65:20:@37541.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 65:20:@37541.4]
  wire  regs_304_io_reset; // @[RegFile.scala 65:20:@37541.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 65:20:@37541.4]
  wire  regs_304_io_enable; // @[RegFile.scala 65:20:@37541.4]
  wire  regs_305_clock; // @[RegFile.scala 65:20:@37555.4]
  wire  regs_305_reset; // @[RegFile.scala 65:20:@37555.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 65:20:@37555.4]
  wire  regs_305_io_reset; // @[RegFile.scala 65:20:@37555.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 65:20:@37555.4]
  wire  regs_305_io_enable; // @[RegFile.scala 65:20:@37555.4]
  wire  regs_306_clock; // @[RegFile.scala 65:20:@37569.4]
  wire  regs_306_reset; // @[RegFile.scala 65:20:@37569.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 65:20:@37569.4]
  wire  regs_306_io_reset; // @[RegFile.scala 65:20:@37569.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 65:20:@37569.4]
  wire  regs_306_io_enable; // @[RegFile.scala 65:20:@37569.4]
  wire  regs_307_clock; // @[RegFile.scala 65:20:@37583.4]
  wire  regs_307_reset; // @[RegFile.scala 65:20:@37583.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 65:20:@37583.4]
  wire  regs_307_io_reset; // @[RegFile.scala 65:20:@37583.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 65:20:@37583.4]
  wire  regs_307_io_enable; // @[RegFile.scala 65:20:@37583.4]
  wire  regs_308_clock; // @[RegFile.scala 65:20:@37597.4]
  wire  regs_308_reset; // @[RegFile.scala 65:20:@37597.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 65:20:@37597.4]
  wire  regs_308_io_reset; // @[RegFile.scala 65:20:@37597.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 65:20:@37597.4]
  wire  regs_308_io_enable; // @[RegFile.scala 65:20:@37597.4]
  wire  regs_309_clock; // @[RegFile.scala 65:20:@37611.4]
  wire  regs_309_reset; // @[RegFile.scala 65:20:@37611.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 65:20:@37611.4]
  wire  regs_309_io_reset; // @[RegFile.scala 65:20:@37611.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 65:20:@37611.4]
  wire  regs_309_io_enable; // @[RegFile.scala 65:20:@37611.4]
  wire  regs_310_clock; // @[RegFile.scala 65:20:@37625.4]
  wire  regs_310_reset; // @[RegFile.scala 65:20:@37625.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 65:20:@37625.4]
  wire  regs_310_io_reset; // @[RegFile.scala 65:20:@37625.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 65:20:@37625.4]
  wire  regs_310_io_enable; // @[RegFile.scala 65:20:@37625.4]
  wire  regs_311_clock; // @[RegFile.scala 65:20:@37639.4]
  wire  regs_311_reset; // @[RegFile.scala 65:20:@37639.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 65:20:@37639.4]
  wire  regs_311_io_reset; // @[RegFile.scala 65:20:@37639.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 65:20:@37639.4]
  wire  regs_311_io_enable; // @[RegFile.scala 65:20:@37639.4]
  wire  regs_312_clock; // @[RegFile.scala 65:20:@37653.4]
  wire  regs_312_reset; // @[RegFile.scala 65:20:@37653.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 65:20:@37653.4]
  wire  regs_312_io_reset; // @[RegFile.scala 65:20:@37653.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 65:20:@37653.4]
  wire  regs_312_io_enable; // @[RegFile.scala 65:20:@37653.4]
  wire  regs_313_clock; // @[RegFile.scala 65:20:@37667.4]
  wire  regs_313_reset; // @[RegFile.scala 65:20:@37667.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 65:20:@37667.4]
  wire  regs_313_io_reset; // @[RegFile.scala 65:20:@37667.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 65:20:@37667.4]
  wire  regs_313_io_enable; // @[RegFile.scala 65:20:@37667.4]
  wire  regs_314_clock; // @[RegFile.scala 65:20:@37681.4]
  wire  regs_314_reset; // @[RegFile.scala 65:20:@37681.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 65:20:@37681.4]
  wire  regs_314_io_reset; // @[RegFile.scala 65:20:@37681.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 65:20:@37681.4]
  wire  regs_314_io_enable; // @[RegFile.scala 65:20:@37681.4]
  wire  regs_315_clock; // @[RegFile.scala 65:20:@37695.4]
  wire  regs_315_reset; // @[RegFile.scala 65:20:@37695.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 65:20:@37695.4]
  wire  regs_315_io_reset; // @[RegFile.scala 65:20:@37695.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 65:20:@37695.4]
  wire  regs_315_io_enable; // @[RegFile.scala 65:20:@37695.4]
  wire  regs_316_clock; // @[RegFile.scala 65:20:@37709.4]
  wire  regs_316_reset; // @[RegFile.scala 65:20:@37709.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 65:20:@37709.4]
  wire  regs_316_io_reset; // @[RegFile.scala 65:20:@37709.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 65:20:@37709.4]
  wire  regs_316_io_enable; // @[RegFile.scala 65:20:@37709.4]
  wire  regs_317_clock; // @[RegFile.scala 65:20:@37723.4]
  wire  regs_317_reset; // @[RegFile.scala 65:20:@37723.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 65:20:@37723.4]
  wire  regs_317_io_reset; // @[RegFile.scala 65:20:@37723.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 65:20:@37723.4]
  wire  regs_317_io_enable; // @[RegFile.scala 65:20:@37723.4]
  wire  regs_318_clock; // @[RegFile.scala 65:20:@37737.4]
  wire  regs_318_reset; // @[RegFile.scala 65:20:@37737.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 65:20:@37737.4]
  wire  regs_318_io_reset; // @[RegFile.scala 65:20:@37737.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 65:20:@37737.4]
  wire  regs_318_io_enable; // @[RegFile.scala 65:20:@37737.4]
  wire  regs_319_clock; // @[RegFile.scala 65:20:@37751.4]
  wire  regs_319_reset; // @[RegFile.scala 65:20:@37751.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 65:20:@37751.4]
  wire  regs_319_io_reset; // @[RegFile.scala 65:20:@37751.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 65:20:@37751.4]
  wire  regs_319_io_enable; // @[RegFile.scala 65:20:@37751.4]
  wire  regs_320_clock; // @[RegFile.scala 65:20:@37765.4]
  wire  regs_320_reset; // @[RegFile.scala 65:20:@37765.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 65:20:@37765.4]
  wire  regs_320_io_reset; // @[RegFile.scala 65:20:@37765.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 65:20:@37765.4]
  wire  regs_320_io_enable; // @[RegFile.scala 65:20:@37765.4]
  wire  regs_321_clock; // @[RegFile.scala 65:20:@37779.4]
  wire  regs_321_reset; // @[RegFile.scala 65:20:@37779.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 65:20:@37779.4]
  wire  regs_321_io_reset; // @[RegFile.scala 65:20:@37779.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 65:20:@37779.4]
  wire  regs_321_io_enable; // @[RegFile.scala 65:20:@37779.4]
  wire  regs_322_clock; // @[RegFile.scala 65:20:@37793.4]
  wire  regs_322_reset; // @[RegFile.scala 65:20:@37793.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 65:20:@37793.4]
  wire  regs_322_io_reset; // @[RegFile.scala 65:20:@37793.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 65:20:@37793.4]
  wire  regs_322_io_enable; // @[RegFile.scala 65:20:@37793.4]
  wire  regs_323_clock; // @[RegFile.scala 65:20:@37807.4]
  wire  regs_323_reset; // @[RegFile.scala 65:20:@37807.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 65:20:@37807.4]
  wire  regs_323_io_reset; // @[RegFile.scala 65:20:@37807.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 65:20:@37807.4]
  wire  regs_323_io_enable; // @[RegFile.scala 65:20:@37807.4]
  wire  regs_324_clock; // @[RegFile.scala 65:20:@37821.4]
  wire  regs_324_reset; // @[RegFile.scala 65:20:@37821.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 65:20:@37821.4]
  wire  regs_324_io_reset; // @[RegFile.scala 65:20:@37821.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 65:20:@37821.4]
  wire  regs_324_io_enable; // @[RegFile.scala 65:20:@37821.4]
  wire  regs_325_clock; // @[RegFile.scala 65:20:@37835.4]
  wire  regs_325_reset; // @[RegFile.scala 65:20:@37835.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 65:20:@37835.4]
  wire  regs_325_io_reset; // @[RegFile.scala 65:20:@37835.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 65:20:@37835.4]
  wire  regs_325_io_enable; // @[RegFile.scala 65:20:@37835.4]
  wire  regs_326_clock; // @[RegFile.scala 65:20:@37849.4]
  wire  regs_326_reset; // @[RegFile.scala 65:20:@37849.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 65:20:@37849.4]
  wire  regs_326_io_reset; // @[RegFile.scala 65:20:@37849.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 65:20:@37849.4]
  wire  regs_326_io_enable; // @[RegFile.scala 65:20:@37849.4]
  wire  regs_327_clock; // @[RegFile.scala 65:20:@37863.4]
  wire  regs_327_reset; // @[RegFile.scala 65:20:@37863.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 65:20:@37863.4]
  wire  regs_327_io_reset; // @[RegFile.scala 65:20:@37863.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 65:20:@37863.4]
  wire  regs_327_io_enable; // @[RegFile.scala 65:20:@37863.4]
  wire  regs_328_clock; // @[RegFile.scala 65:20:@37877.4]
  wire  regs_328_reset; // @[RegFile.scala 65:20:@37877.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 65:20:@37877.4]
  wire  regs_328_io_reset; // @[RegFile.scala 65:20:@37877.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 65:20:@37877.4]
  wire  regs_328_io_enable; // @[RegFile.scala 65:20:@37877.4]
  wire  regs_329_clock; // @[RegFile.scala 65:20:@37891.4]
  wire  regs_329_reset; // @[RegFile.scala 65:20:@37891.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 65:20:@37891.4]
  wire  regs_329_io_reset; // @[RegFile.scala 65:20:@37891.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 65:20:@37891.4]
  wire  regs_329_io_enable; // @[RegFile.scala 65:20:@37891.4]
  wire  regs_330_clock; // @[RegFile.scala 65:20:@37905.4]
  wire  regs_330_reset; // @[RegFile.scala 65:20:@37905.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 65:20:@37905.4]
  wire  regs_330_io_reset; // @[RegFile.scala 65:20:@37905.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 65:20:@37905.4]
  wire  regs_330_io_enable; // @[RegFile.scala 65:20:@37905.4]
  wire  regs_331_clock; // @[RegFile.scala 65:20:@37919.4]
  wire  regs_331_reset; // @[RegFile.scala 65:20:@37919.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 65:20:@37919.4]
  wire  regs_331_io_reset; // @[RegFile.scala 65:20:@37919.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 65:20:@37919.4]
  wire  regs_331_io_enable; // @[RegFile.scala 65:20:@37919.4]
  wire  regs_332_clock; // @[RegFile.scala 65:20:@37933.4]
  wire  regs_332_reset; // @[RegFile.scala 65:20:@37933.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 65:20:@37933.4]
  wire  regs_332_io_reset; // @[RegFile.scala 65:20:@37933.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 65:20:@37933.4]
  wire  regs_332_io_enable; // @[RegFile.scala 65:20:@37933.4]
  wire  regs_333_clock; // @[RegFile.scala 65:20:@37947.4]
  wire  regs_333_reset; // @[RegFile.scala 65:20:@37947.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 65:20:@37947.4]
  wire  regs_333_io_reset; // @[RegFile.scala 65:20:@37947.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 65:20:@37947.4]
  wire  regs_333_io_enable; // @[RegFile.scala 65:20:@37947.4]
  wire  regs_334_clock; // @[RegFile.scala 65:20:@37961.4]
  wire  regs_334_reset; // @[RegFile.scala 65:20:@37961.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 65:20:@37961.4]
  wire  regs_334_io_reset; // @[RegFile.scala 65:20:@37961.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 65:20:@37961.4]
  wire  regs_334_io_enable; // @[RegFile.scala 65:20:@37961.4]
  wire  regs_335_clock; // @[RegFile.scala 65:20:@37975.4]
  wire  regs_335_reset; // @[RegFile.scala 65:20:@37975.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 65:20:@37975.4]
  wire  regs_335_io_reset; // @[RegFile.scala 65:20:@37975.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 65:20:@37975.4]
  wire  regs_335_io_enable; // @[RegFile.scala 65:20:@37975.4]
  wire  regs_336_clock; // @[RegFile.scala 65:20:@37989.4]
  wire  regs_336_reset; // @[RegFile.scala 65:20:@37989.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 65:20:@37989.4]
  wire  regs_336_io_reset; // @[RegFile.scala 65:20:@37989.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 65:20:@37989.4]
  wire  regs_336_io_enable; // @[RegFile.scala 65:20:@37989.4]
  wire  regs_337_clock; // @[RegFile.scala 65:20:@38003.4]
  wire  regs_337_reset; // @[RegFile.scala 65:20:@38003.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 65:20:@38003.4]
  wire  regs_337_io_reset; // @[RegFile.scala 65:20:@38003.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 65:20:@38003.4]
  wire  regs_337_io_enable; // @[RegFile.scala 65:20:@38003.4]
  wire  regs_338_clock; // @[RegFile.scala 65:20:@38017.4]
  wire  regs_338_reset; // @[RegFile.scala 65:20:@38017.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 65:20:@38017.4]
  wire  regs_338_io_reset; // @[RegFile.scala 65:20:@38017.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 65:20:@38017.4]
  wire  regs_338_io_enable; // @[RegFile.scala 65:20:@38017.4]
  wire  regs_339_clock; // @[RegFile.scala 65:20:@38031.4]
  wire  regs_339_reset; // @[RegFile.scala 65:20:@38031.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 65:20:@38031.4]
  wire  regs_339_io_reset; // @[RegFile.scala 65:20:@38031.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 65:20:@38031.4]
  wire  regs_339_io_enable; // @[RegFile.scala 65:20:@38031.4]
  wire  regs_340_clock; // @[RegFile.scala 65:20:@38045.4]
  wire  regs_340_reset; // @[RegFile.scala 65:20:@38045.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 65:20:@38045.4]
  wire  regs_340_io_reset; // @[RegFile.scala 65:20:@38045.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 65:20:@38045.4]
  wire  regs_340_io_enable; // @[RegFile.scala 65:20:@38045.4]
  wire  regs_341_clock; // @[RegFile.scala 65:20:@38059.4]
  wire  regs_341_reset; // @[RegFile.scala 65:20:@38059.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 65:20:@38059.4]
  wire  regs_341_io_reset; // @[RegFile.scala 65:20:@38059.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 65:20:@38059.4]
  wire  regs_341_io_enable; // @[RegFile.scala 65:20:@38059.4]
  wire  regs_342_clock; // @[RegFile.scala 65:20:@38073.4]
  wire  regs_342_reset; // @[RegFile.scala 65:20:@38073.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 65:20:@38073.4]
  wire  regs_342_io_reset; // @[RegFile.scala 65:20:@38073.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 65:20:@38073.4]
  wire  regs_342_io_enable; // @[RegFile.scala 65:20:@38073.4]
  wire  regs_343_clock; // @[RegFile.scala 65:20:@38087.4]
  wire  regs_343_reset; // @[RegFile.scala 65:20:@38087.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 65:20:@38087.4]
  wire  regs_343_io_reset; // @[RegFile.scala 65:20:@38087.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 65:20:@38087.4]
  wire  regs_343_io_enable; // @[RegFile.scala 65:20:@38087.4]
  wire  regs_344_clock; // @[RegFile.scala 65:20:@38101.4]
  wire  regs_344_reset; // @[RegFile.scala 65:20:@38101.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 65:20:@38101.4]
  wire  regs_344_io_reset; // @[RegFile.scala 65:20:@38101.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 65:20:@38101.4]
  wire  regs_344_io_enable; // @[RegFile.scala 65:20:@38101.4]
  wire  regs_345_clock; // @[RegFile.scala 65:20:@38115.4]
  wire  regs_345_reset; // @[RegFile.scala 65:20:@38115.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 65:20:@38115.4]
  wire  regs_345_io_reset; // @[RegFile.scala 65:20:@38115.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 65:20:@38115.4]
  wire  regs_345_io_enable; // @[RegFile.scala 65:20:@38115.4]
  wire  regs_346_clock; // @[RegFile.scala 65:20:@38129.4]
  wire  regs_346_reset; // @[RegFile.scala 65:20:@38129.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 65:20:@38129.4]
  wire  regs_346_io_reset; // @[RegFile.scala 65:20:@38129.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 65:20:@38129.4]
  wire  regs_346_io_enable; // @[RegFile.scala 65:20:@38129.4]
  wire  regs_347_clock; // @[RegFile.scala 65:20:@38143.4]
  wire  regs_347_reset; // @[RegFile.scala 65:20:@38143.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 65:20:@38143.4]
  wire  regs_347_io_reset; // @[RegFile.scala 65:20:@38143.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 65:20:@38143.4]
  wire  regs_347_io_enable; // @[RegFile.scala 65:20:@38143.4]
  wire  regs_348_clock; // @[RegFile.scala 65:20:@38157.4]
  wire  regs_348_reset; // @[RegFile.scala 65:20:@38157.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 65:20:@38157.4]
  wire  regs_348_io_reset; // @[RegFile.scala 65:20:@38157.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 65:20:@38157.4]
  wire  regs_348_io_enable; // @[RegFile.scala 65:20:@38157.4]
  wire  regs_349_clock; // @[RegFile.scala 65:20:@38171.4]
  wire  regs_349_reset; // @[RegFile.scala 65:20:@38171.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 65:20:@38171.4]
  wire  regs_349_io_reset; // @[RegFile.scala 65:20:@38171.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 65:20:@38171.4]
  wire  regs_349_io_enable; // @[RegFile.scala 65:20:@38171.4]
  wire  regs_350_clock; // @[RegFile.scala 65:20:@38185.4]
  wire  regs_350_reset; // @[RegFile.scala 65:20:@38185.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 65:20:@38185.4]
  wire  regs_350_io_reset; // @[RegFile.scala 65:20:@38185.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 65:20:@38185.4]
  wire  regs_350_io_enable; // @[RegFile.scala 65:20:@38185.4]
  wire  regs_351_clock; // @[RegFile.scala 65:20:@38199.4]
  wire  regs_351_reset; // @[RegFile.scala 65:20:@38199.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 65:20:@38199.4]
  wire  regs_351_io_reset; // @[RegFile.scala 65:20:@38199.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 65:20:@38199.4]
  wire  regs_351_io_enable; // @[RegFile.scala 65:20:@38199.4]
  wire  regs_352_clock; // @[RegFile.scala 65:20:@38213.4]
  wire  regs_352_reset; // @[RegFile.scala 65:20:@38213.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 65:20:@38213.4]
  wire  regs_352_io_reset; // @[RegFile.scala 65:20:@38213.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 65:20:@38213.4]
  wire  regs_352_io_enable; // @[RegFile.scala 65:20:@38213.4]
  wire  regs_353_clock; // @[RegFile.scala 65:20:@38227.4]
  wire  regs_353_reset; // @[RegFile.scala 65:20:@38227.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 65:20:@38227.4]
  wire  regs_353_io_reset; // @[RegFile.scala 65:20:@38227.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 65:20:@38227.4]
  wire  regs_353_io_enable; // @[RegFile.scala 65:20:@38227.4]
  wire  regs_354_clock; // @[RegFile.scala 65:20:@38241.4]
  wire  regs_354_reset; // @[RegFile.scala 65:20:@38241.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 65:20:@38241.4]
  wire  regs_354_io_reset; // @[RegFile.scala 65:20:@38241.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 65:20:@38241.4]
  wire  regs_354_io_enable; // @[RegFile.scala 65:20:@38241.4]
  wire  regs_355_clock; // @[RegFile.scala 65:20:@38255.4]
  wire  regs_355_reset; // @[RegFile.scala 65:20:@38255.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 65:20:@38255.4]
  wire  regs_355_io_reset; // @[RegFile.scala 65:20:@38255.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 65:20:@38255.4]
  wire  regs_355_io_enable; // @[RegFile.scala 65:20:@38255.4]
  wire  regs_356_clock; // @[RegFile.scala 65:20:@38269.4]
  wire  regs_356_reset; // @[RegFile.scala 65:20:@38269.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 65:20:@38269.4]
  wire  regs_356_io_reset; // @[RegFile.scala 65:20:@38269.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 65:20:@38269.4]
  wire  regs_356_io_enable; // @[RegFile.scala 65:20:@38269.4]
  wire  regs_357_clock; // @[RegFile.scala 65:20:@38283.4]
  wire  regs_357_reset; // @[RegFile.scala 65:20:@38283.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 65:20:@38283.4]
  wire  regs_357_io_reset; // @[RegFile.scala 65:20:@38283.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 65:20:@38283.4]
  wire  regs_357_io_enable; // @[RegFile.scala 65:20:@38283.4]
  wire  regs_358_clock; // @[RegFile.scala 65:20:@38297.4]
  wire  regs_358_reset; // @[RegFile.scala 65:20:@38297.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 65:20:@38297.4]
  wire  regs_358_io_reset; // @[RegFile.scala 65:20:@38297.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 65:20:@38297.4]
  wire  regs_358_io_enable; // @[RegFile.scala 65:20:@38297.4]
  wire  regs_359_clock; // @[RegFile.scala 65:20:@38311.4]
  wire  regs_359_reset; // @[RegFile.scala 65:20:@38311.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 65:20:@38311.4]
  wire  regs_359_io_reset; // @[RegFile.scala 65:20:@38311.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 65:20:@38311.4]
  wire  regs_359_io_enable; // @[RegFile.scala 65:20:@38311.4]
  wire  regs_360_clock; // @[RegFile.scala 65:20:@38325.4]
  wire  regs_360_reset; // @[RegFile.scala 65:20:@38325.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 65:20:@38325.4]
  wire  regs_360_io_reset; // @[RegFile.scala 65:20:@38325.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 65:20:@38325.4]
  wire  regs_360_io_enable; // @[RegFile.scala 65:20:@38325.4]
  wire  regs_361_clock; // @[RegFile.scala 65:20:@38339.4]
  wire  regs_361_reset; // @[RegFile.scala 65:20:@38339.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 65:20:@38339.4]
  wire  regs_361_io_reset; // @[RegFile.scala 65:20:@38339.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 65:20:@38339.4]
  wire  regs_361_io_enable; // @[RegFile.scala 65:20:@38339.4]
  wire  regs_362_clock; // @[RegFile.scala 65:20:@38353.4]
  wire  regs_362_reset; // @[RegFile.scala 65:20:@38353.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 65:20:@38353.4]
  wire  regs_362_io_reset; // @[RegFile.scala 65:20:@38353.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 65:20:@38353.4]
  wire  regs_362_io_enable; // @[RegFile.scala 65:20:@38353.4]
  wire  regs_363_clock; // @[RegFile.scala 65:20:@38367.4]
  wire  regs_363_reset; // @[RegFile.scala 65:20:@38367.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 65:20:@38367.4]
  wire  regs_363_io_reset; // @[RegFile.scala 65:20:@38367.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 65:20:@38367.4]
  wire  regs_363_io_enable; // @[RegFile.scala 65:20:@38367.4]
  wire  regs_364_clock; // @[RegFile.scala 65:20:@38381.4]
  wire  regs_364_reset; // @[RegFile.scala 65:20:@38381.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 65:20:@38381.4]
  wire  regs_364_io_reset; // @[RegFile.scala 65:20:@38381.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 65:20:@38381.4]
  wire  regs_364_io_enable; // @[RegFile.scala 65:20:@38381.4]
  wire  regs_365_clock; // @[RegFile.scala 65:20:@38395.4]
  wire  regs_365_reset; // @[RegFile.scala 65:20:@38395.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 65:20:@38395.4]
  wire  regs_365_io_reset; // @[RegFile.scala 65:20:@38395.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 65:20:@38395.4]
  wire  regs_365_io_enable; // @[RegFile.scala 65:20:@38395.4]
  wire  regs_366_clock; // @[RegFile.scala 65:20:@38409.4]
  wire  regs_366_reset; // @[RegFile.scala 65:20:@38409.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 65:20:@38409.4]
  wire  regs_366_io_reset; // @[RegFile.scala 65:20:@38409.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 65:20:@38409.4]
  wire  regs_366_io_enable; // @[RegFile.scala 65:20:@38409.4]
  wire  regs_367_clock; // @[RegFile.scala 65:20:@38423.4]
  wire  regs_367_reset; // @[RegFile.scala 65:20:@38423.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 65:20:@38423.4]
  wire  regs_367_io_reset; // @[RegFile.scala 65:20:@38423.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 65:20:@38423.4]
  wire  regs_367_io_enable; // @[RegFile.scala 65:20:@38423.4]
  wire  regs_368_clock; // @[RegFile.scala 65:20:@38437.4]
  wire  regs_368_reset; // @[RegFile.scala 65:20:@38437.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 65:20:@38437.4]
  wire  regs_368_io_reset; // @[RegFile.scala 65:20:@38437.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 65:20:@38437.4]
  wire  regs_368_io_enable; // @[RegFile.scala 65:20:@38437.4]
  wire  regs_369_clock; // @[RegFile.scala 65:20:@38451.4]
  wire  regs_369_reset; // @[RegFile.scala 65:20:@38451.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 65:20:@38451.4]
  wire  regs_369_io_reset; // @[RegFile.scala 65:20:@38451.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 65:20:@38451.4]
  wire  regs_369_io_enable; // @[RegFile.scala 65:20:@38451.4]
  wire  regs_370_clock; // @[RegFile.scala 65:20:@38465.4]
  wire  regs_370_reset; // @[RegFile.scala 65:20:@38465.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 65:20:@38465.4]
  wire  regs_370_io_reset; // @[RegFile.scala 65:20:@38465.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 65:20:@38465.4]
  wire  regs_370_io_enable; // @[RegFile.scala 65:20:@38465.4]
  wire  regs_371_clock; // @[RegFile.scala 65:20:@38479.4]
  wire  regs_371_reset; // @[RegFile.scala 65:20:@38479.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 65:20:@38479.4]
  wire  regs_371_io_reset; // @[RegFile.scala 65:20:@38479.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 65:20:@38479.4]
  wire  regs_371_io_enable; // @[RegFile.scala 65:20:@38479.4]
  wire  regs_372_clock; // @[RegFile.scala 65:20:@38493.4]
  wire  regs_372_reset; // @[RegFile.scala 65:20:@38493.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 65:20:@38493.4]
  wire  regs_372_io_reset; // @[RegFile.scala 65:20:@38493.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 65:20:@38493.4]
  wire  regs_372_io_enable; // @[RegFile.scala 65:20:@38493.4]
  wire  regs_373_clock; // @[RegFile.scala 65:20:@38507.4]
  wire  regs_373_reset; // @[RegFile.scala 65:20:@38507.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 65:20:@38507.4]
  wire  regs_373_io_reset; // @[RegFile.scala 65:20:@38507.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 65:20:@38507.4]
  wire  regs_373_io_enable; // @[RegFile.scala 65:20:@38507.4]
  wire  regs_374_clock; // @[RegFile.scala 65:20:@38521.4]
  wire  regs_374_reset; // @[RegFile.scala 65:20:@38521.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 65:20:@38521.4]
  wire  regs_374_io_reset; // @[RegFile.scala 65:20:@38521.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 65:20:@38521.4]
  wire  regs_374_io_enable; // @[RegFile.scala 65:20:@38521.4]
  wire  regs_375_clock; // @[RegFile.scala 65:20:@38535.4]
  wire  regs_375_reset; // @[RegFile.scala 65:20:@38535.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 65:20:@38535.4]
  wire  regs_375_io_reset; // @[RegFile.scala 65:20:@38535.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 65:20:@38535.4]
  wire  regs_375_io_enable; // @[RegFile.scala 65:20:@38535.4]
  wire  regs_376_clock; // @[RegFile.scala 65:20:@38549.4]
  wire  regs_376_reset; // @[RegFile.scala 65:20:@38549.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 65:20:@38549.4]
  wire  regs_376_io_reset; // @[RegFile.scala 65:20:@38549.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 65:20:@38549.4]
  wire  regs_376_io_enable; // @[RegFile.scala 65:20:@38549.4]
  wire  regs_377_clock; // @[RegFile.scala 65:20:@38563.4]
  wire  regs_377_reset; // @[RegFile.scala 65:20:@38563.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 65:20:@38563.4]
  wire  regs_377_io_reset; // @[RegFile.scala 65:20:@38563.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 65:20:@38563.4]
  wire  regs_377_io_enable; // @[RegFile.scala 65:20:@38563.4]
  wire  regs_378_clock; // @[RegFile.scala 65:20:@38577.4]
  wire  regs_378_reset; // @[RegFile.scala 65:20:@38577.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 65:20:@38577.4]
  wire  regs_378_io_reset; // @[RegFile.scala 65:20:@38577.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 65:20:@38577.4]
  wire  regs_378_io_enable; // @[RegFile.scala 65:20:@38577.4]
  wire  regs_379_clock; // @[RegFile.scala 65:20:@38591.4]
  wire  regs_379_reset; // @[RegFile.scala 65:20:@38591.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 65:20:@38591.4]
  wire  regs_379_io_reset; // @[RegFile.scala 65:20:@38591.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 65:20:@38591.4]
  wire  regs_379_io_enable; // @[RegFile.scala 65:20:@38591.4]
  wire  regs_380_clock; // @[RegFile.scala 65:20:@38605.4]
  wire  regs_380_reset; // @[RegFile.scala 65:20:@38605.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 65:20:@38605.4]
  wire  regs_380_io_reset; // @[RegFile.scala 65:20:@38605.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 65:20:@38605.4]
  wire  regs_380_io_enable; // @[RegFile.scala 65:20:@38605.4]
  wire  regs_381_clock; // @[RegFile.scala 65:20:@38619.4]
  wire  regs_381_reset; // @[RegFile.scala 65:20:@38619.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 65:20:@38619.4]
  wire  regs_381_io_reset; // @[RegFile.scala 65:20:@38619.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 65:20:@38619.4]
  wire  regs_381_io_enable; // @[RegFile.scala 65:20:@38619.4]
  wire  regs_382_clock; // @[RegFile.scala 65:20:@38633.4]
  wire  regs_382_reset; // @[RegFile.scala 65:20:@38633.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 65:20:@38633.4]
  wire  regs_382_io_reset; // @[RegFile.scala 65:20:@38633.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 65:20:@38633.4]
  wire  regs_382_io_enable; // @[RegFile.scala 65:20:@38633.4]
  wire  regs_383_clock; // @[RegFile.scala 65:20:@38647.4]
  wire  regs_383_reset; // @[RegFile.scala 65:20:@38647.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 65:20:@38647.4]
  wire  regs_383_io_reset; // @[RegFile.scala 65:20:@38647.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 65:20:@38647.4]
  wire  regs_383_io_enable; // @[RegFile.scala 65:20:@38647.4]
  wire  regs_384_clock; // @[RegFile.scala 65:20:@38661.4]
  wire  regs_384_reset; // @[RegFile.scala 65:20:@38661.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 65:20:@38661.4]
  wire  regs_384_io_reset; // @[RegFile.scala 65:20:@38661.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 65:20:@38661.4]
  wire  regs_384_io_enable; // @[RegFile.scala 65:20:@38661.4]
  wire  regs_385_clock; // @[RegFile.scala 65:20:@38675.4]
  wire  regs_385_reset; // @[RegFile.scala 65:20:@38675.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 65:20:@38675.4]
  wire  regs_385_io_reset; // @[RegFile.scala 65:20:@38675.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 65:20:@38675.4]
  wire  regs_385_io_enable; // @[RegFile.scala 65:20:@38675.4]
  wire  regs_386_clock; // @[RegFile.scala 65:20:@38689.4]
  wire  regs_386_reset; // @[RegFile.scala 65:20:@38689.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 65:20:@38689.4]
  wire  regs_386_io_reset; // @[RegFile.scala 65:20:@38689.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 65:20:@38689.4]
  wire  regs_386_io_enable; // @[RegFile.scala 65:20:@38689.4]
  wire  regs_387_clock; // @[RegFile.scala 65:20:@38703.4]
  wire  regs_387_reset; // @[RegFile.scala 65:20:@38703.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 65:20:@38703.4]
  wire  regs_387_io_reset; // @[RegFile.scala 65:20:@38703.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 65:20:@38703.4]
  wire  regs_387_io_enable; // @[RegFile.scala 65:20:@38703.4]
  wire  regs_388_clock; // @[RegFile.scala 65:20:@38717.4]
  wire  regs_388_reset; // @[RegFile.scala 65:20:@38717.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 65:20:@38717.4]
  wire  regs_388_io_reset; // @[RegFile.scala 65:20:@38717.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 65:20:@38717.4]
  wire  regs_388_io_enable; // @[RegFile.scala 65:20:@38717.4]
  wire  regs_389_clock; // @[RegFile.scala 65:20:@38731.4]
  wire  regs_389_reset; // @[RegFile.scala 65:20:@38731.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 65:20:@38731.4]
  wire  regs_389_io_reset; // @[RegFile.scala 65:20:@38731.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 65:20:@38731.4]
  wire  regs_389_io_enable; // @[RegFile.scala 65:20:@38731.4]
  wire  regs_390_clock; // @[RegFile.scala 65:20:@38745.4]
  wire  regs_390_reset; // @[RegFile.scala 65:20:@38745.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 65:20:@38745.4]
  wire  regs_390_io_reset; // @[RegFile.scala 65:20:@38745.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 65:20:@38745.4]
  wire  regs_390_io_enable; // @[RegFile.scala 65:20:@38745.4]
  wire  regs_391_clock; // @[RegFile.scala 65:20:@38759.4]
  wire  regs_391_reset; // @[RegFile.scala 65:20:@38759.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 65:20:@38759.4]
  wire  regs_391_io_reset; // @[RegFile.scala 65:20:@38759.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 65:20:@38759.4]
  wire  regs_391_io_enable; // @[RegFile.scala 65:20:@38759.4]
  wire  regs_392_clock; // @[RegFile.scala 65:20:@38773.4]
  wire  regs_392_reset; // @[RegFile.scala 65:20:@38773.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 65:20:@38773.4]
  wire  regs_392_io_reset; // @[RegFile.scala 65:20:@38773.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 65:20:@38773.4]
  wire  regs_392_io_enable; // @[RegFile.scala 65:20:@38773.4]
  wire  regs_393_clock; // @[RegFile.scala 65:20:@38787.4]
  wire  regs_393_reset; // @[RegFile.scala 65:20:@38787.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 65:20:@38787.4]
  wire  regs_393_io_reset; // @[RegFile.scala 65:20:@38787.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 65:20:@38787.4]
  wire  regs_393_io_enable; // @[RegFile.scala 65:20:@38787.4]
  wire  regs_394_clock; // @[RegFile.scala 65:20:@38801.4]
  wire  regs_394_reset; // @[RegFile.scala 65:20:@38801.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 65:20:@38801.4]
  wire  regs_394_io_reset; // @[RegFile.scala 65:20:@38801.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 65:20:@38801.4]
  wire  regs_394_io_enable; // @[RegFile.scala 65:20:@38801.4]
  wire  regs_395_clock; // @[RegFile.scala 65:20:@38815.4]
  wire  regs_395_reset; // @[RegFile.scala 65:20:@38815.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 65:20:@38815.4]
  wire  regs_395_io_reset; // @[RegFile.scala 65:20:@38815.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 65:20:@38815.4]
  wire  regs_395_io_enable; // @[RegFile.scala 65:20:@38815.4]
  wire  regs_396_clock; // @[RegFile.scala 65:20:@38829.4]
  wire  regs_396_reset; // @[RegFile.scala 65:20:@38829.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 65:20:@38829.4]
  wire  regs_396_io_reset; // @[RegFile.scala 65:20:@38829.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 65:20:@38829.4]
  wire  regs_396_io_enable; // @[RegFile.scala 65:20:@38829.4]
  wire  regs_397_clock; // @[RegFile.scala 65:20:@38843.4]
  wire  regs_397_reset; // @[RegFile.scala 65:20:@38843.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 65:20:@38843.4]
  wire  regs_397_io_reset; // @[RegFile.scala 65:20:@38843.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 65:20:@38843.4]
  wire  regs_397_io_enable; // @[RegFile.scala 65:20:@38843.4]
  wire  regs_398_clock; // @[RegFile.scala 65:20:@38857.4]
  wire  regs_398_reset; // @[RegFile.scala 65:20:@38857.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 65:20:@38857.4]
  wire  regs_398_io_reset; // @[RegFile.scala 65:20:@38857.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 65:20:@38857.4]
  wire  regs_398_io_enable; // @[RegFile.scala 65:20:@38857.4]
  wire  regs_399_clock; // @[RegFile.scala 65:20:@38871.4]
  wire  regs_399_reset; // @[RegFile.scala 65:20:@38871.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 65:20:@38871.4]
  wire  regs_399_io_reset; // @[RegFile.scala 65:20:@38871.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 65:20:@38871.4]
  wire  regs_399_io_enable; // @[RegFile.scala 65:20:@38871.4]
  wire  regs_400_clock; // @[RegFile.scala 65:20:@38885.4]
  wire  regs_400_reset; // @[RegFile.scala 65:20:@38885.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 65:20:@38885.4]
  wire  regs_400_io_reset; // @[RegFile.scala 65:20:@38885.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 65:20:@38885.4]
  wire  regs_400_io_enable; // @[RegFile.scala 65:20:@38885.4]
  wire  regs_401_clock; // @[RegFile.scala 65:20:@38899.4]
  wire  regs_401_reset; // @[RegFile.scala 65:20:@38899.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 65:20:@38899.4]
  wire  regs_401_io_reset; // @[RegFile.scala 65:20:@38899.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 65:20:@38899.4]
  wire  regs_401_io_enable; // @[RegFile.scala 65:20:@38899.4]
  wire  regs_402_clock; // @[RegFile.scala 65:20:@38913.4]
  wire  regs_402_reset; // @[RegFile.scala 65:20:@38913.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 65:20:@38913.4]
  wire  regs_402_io_reset; // @[RegFile.scala 65:20:@38913.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 65:20:@38913.4]
  wire  regs_402_io_enable; // @[RegFile.scala 65:20:@38913.4]
  wire  regs_403_clock; // @[RegFile.scala 65:20:@38927.4]
  wire  regs_403_reset; // @[RegFile.scala 65:20:@38927.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 65:20:@38927.4]
  wire  regs_403_io_reset; // @[RegFile.scala 65:20:@38927.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 65:20:@38927.4]
  wire  regs_403_io_enable; // @[RegFile.scala 65:20:@38927.4]
  wire  regs_404_clock; // @[RegFile.scala 65:20:@38941.4]
  wire  regs_404_reset; // @[RegFile.scala 65:20:@38941.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 65:20:@38941.4]
  wire  regs_404_io_reset; // @[RegFile.scala 65:20:@38941.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 65:20:@38941.4]
  wire  regs_404_io_enable; // @[RegFile.scala 65:20:@38941.4]
  wire  regs_405_clock; // @[RegFile.scala 65:20:@38955.4]
  wire  regs_405_reset; // @[RegFile.scala 65:20:@38955.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 65:20:@38955.4]
  wire  regs_405_io_reset; // @[RegFile.scala 65:20:@38955.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 65:20:@38955.4]
  wire  regs_405_io_enable; // @[RegFile.scala 65:20:@38955.4]
  wire  regs_406_clock; // @[RegFile.scala 65:20:@38969.4]
  wire  regs_406_reset; // @[RegFile.scala 65:20:@38969.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 65:20:@38969.4]
  wire  regs_406_io_reset; // @[RegFile.scala 65:20:@38969.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 65:20:@38969.4]
  wire  regs_406_io_enable; // @[RegFile.scala 65:20:@38969.4]
  wire  regs_407_clock; // @[RegFile.scala 65:20:@38983.4]
  wire  regs_407_reset; // @[RegFile.scala 65:20:@38983.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 65:20:@38983.4]
  wire  regs_407_io_reset; // @[RegFile.scala 65:20:@38983.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 65:20:@38983.4]
  wire  regs_407_io_enable; // @[RegFile.scala 65:20:@38983.4]
  wire  regs_408_clock; // @[RegFile.scala 65:20:@38997.4]
  wire  regs_408_reset; // @[RegFile.scala 65:20:@38997.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 65:20:@38997.4]
  wire  regs_408_io_reset; // @[RegFile.scala 65:20:@38997.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 65:20:@38997.4]
  wire  regs_408_io_enable; // @[RegFile.scala 65:20:@38997.4]
  wire  regs_409_clock; // @[RegFile.scala 65:20:@39011.4]
  wire  regs_409_reset; // @[RegFile.scala 65:20:@39011.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 65:20:@39011.4]
  wire  regs_409_io_reset; // @[RegFile.scala 65:20:@39011.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 65:20:@39011.4]
  wire  regs_409_io_enable; // @[RegFile.scala 65:20:@39011.4]
  wire  regs_410_clock; // @[RegFile.scala 65:20:@39025.4]
  wire  regs_410_reset; // @[RegFile.scala 65:20:@39025.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 65:20:@39025.4]
  wire  regs_410_io_reset; // @[RegFile.scala 65:20:@39025.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 65:20:@39025.4]
  wire  regs_410_io_enable; // @[RegFile.scala 65:20:@39025.4]
  wire  regs_411_clock; // @[RegFile.scala 65:20:@39039.4]
  wire  regs_411_reset; // @[RegFile.scala 65:20:@39039.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 65:20:@39039.4]
  wire  regs_411_io_reset; // @[RegFile.scala 65:20:@39039.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 65:20:@39039.4]
  wire  regs_411_io_enable; // @[RegFile.scala 65:20:@39039.4]
  wire  regs_412_clock; // @[RegFile.scala 65:20:@39053.4]
  wire  regs_412_reset; // @[RegFile.scala 65:20:@39053.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 65:20:@39053.4]
  wire  regs_412_io_reset; // @[RegFile.scala 65:20:@39053.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 65:20:@39053.4]
  wire  regs_412_io_enable; // @[RegFile.scala 65:20:@39053.4]
  wire  regs_413_clock; // @[RegFile.scala 65:20:@39067.4]
  wire  regs_413_reset; // @[RegFile.scala 65:20:@39067.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 65:20:@39067.4]
  wire  regs_413_io_reset; // @[RegFile.scala 65:20:@39067.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 65:20:@39067.4]
  wire  regs_413_io_enable; // @[RegFile.scala 65:20:@39067.4]
  wire  regs_414_clock; // @[RegFile.scala 65:20:@39081.4]
  wire  regs_414_reset; // @[RegFile.scala 65:20:@39081.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 65:20:@39081.4]
  wire  regs_414_io_reset; // @[RegFile.scala 65:20:@39081.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 65:20:@39081.4]
  wire  regs_414_io_enable; // @[RegFile.scala 65:20:@39081.4]
  wire  regs_415_clock; // @[RegFile.scala 65:20:@39095.4]
  wire  regs_415_reset; // @[RegFile.scala 65:20:@39095.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 65:20:@39095.4]
  wire  regs_415_io_reset; // @[RegFile.scala 65:20:@39095.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 65:20:@39095.4]
  wire  regs_415_io_enable; // @[RegFile.scala 65:20:@39095.4]
  wire  regs_416_clock; // @[RegFile.scala 65:20:@39109.4]
  wire  regs_416_reset; // @[RegFile.scala 65:20:@39109.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 65:20:@39109.4]
  wire  regs_416_io_reset; // @[RegFile.scala 65:20:@39109.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 65:20:@39109.4]
  wire  regs_416_io_enable; // @[RegFile.scala 65:20:@39109.4]
  wire  regs_417_clock; // @[RegFile.scala 65:20:@39123.4]
  wire  regs_417_reset; // @[RegFile.scala 65:20:@39123.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 65:20:@39123.4]
  wire  regs_417_io_reset; // @[RegFile.scala 65:20:@39123.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 65:20:@39123.4]
  wire  regs_417_io_enable; // @[RegFile.scala 65:20:@39123.4]
  wire  regs_418_clock; // @[RegFile.scala 65:20:@39137.4]
  wire  regs_418_reset; // @[RegFile.scala 65:20:@39137.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 65:20:@39137.4]
  wire  regs_418_io_reset; // @[RegFile.scala 65:20:@39137.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 65:20:@39137.4]
  wire  regs_418_io_enable; // @[RegFile.scala 65:20:@39137.4]
  wire  regs_419_clock; // @[RegFile.scala 65:20:@39151.4]
  wire  regs_419_reset; // @[RegFile.scala 65:20:@39151.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 65:20:@39151.4]
  wire  regs_419_io_reset; // @[RegFile.scala 65:20:@39151.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 65:20:@39151.4]
  wire  regs_419_io_enable; // @[RegFile.scala 65:20:@39151.4]
  wire  regs_420_clock; // @[RegFile.scala 65:20:@39165.4]
  wire  regs_420_reset; // @[RegFile.scala 65:20:@39165.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 65:20:@39165.4]
  wire  regs_420_io_reset; // @[RegFile.scala 65:20:@39165.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 65:20:@39165.4]
  wire  regs_420_io_enable; // @[RegFile.scala 65:20:@39165.4]
  wire  regs_421_clock; // @[RegFile.scala 65:20:@39179.4]
  wire  regs_421_reset; // @[RegFile.scala 65:20:@39179.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 65:20:@39179.4]
  wire  regs_421_io_reset; // @[RegFile.scala 65:20:@39179.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 65:20:@39179.4]
  wire  regs_421_io_enable; // @[RegFile.scala 65:20:@39179.4]
  wire  regs_422_clock; // @[RegFile.scala 65:20:@39193.4]
  wire  regs_422_reset; // @[RegFile.scala 65:20:@39193.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 65:20:@39193.4]
  wire  regs_422_io_reset; // @[RegFile.scala 65:20:@39193.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 65:20:@39193.4]
  wire  regs_422_io_enable; // @[RegFile.scala 65:20:@39193.4]
  wire  regs_423_clock; // @[RegFile.scala 65:20:@39207.4]
  wire  regs_423_reset; // @[RegFile.scala 65:20:@39207.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 65:20:@39207.4]
  wire  regs_423_io_reset; // @[RegFile.scala 65:20:@39207.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 65:20:@39207.4]
  wire  regs_423_io_enable; // @[RegFile.scala 65:20:@39207.4]
  wire  regs_424_clock; // @[RegFile.scala 65:20:@39221.4]
  wire  regs_424_reset; // @[RegFile.scala 65:20:@39221.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 65:20:@39221.4]
  wire  regs_424_io_reset; // @[RegFile.scala 65:20:@39221.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 65:20:@39221.4]
  wire  regs_424_io_enable; // @[RegFile.scala 65:20:@39221.4]
  wire  regs_425_clock; // @[RegFile.scala 65:20:@39235.4]
  wire  regs_425_reset; // @[RegFile.scala 65:20:@39235.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 65:20:@39235.4]
  wire  regs_425_io_reset; // @[RegFile.scala 65:20:@39235.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 65:20:@39235.4]
  wire  regs_425_io_enable; // @[RegFile.scala 65:20:@39235.4]
  wire  regs_426_clock; // @[RegFile.scala 65:20:@39249.4]
  wire  regs_426_reset; // @[RegFile.scala 65:20:@39249.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 65:20:@39249.4]
  wire  regs_426_io_reset; // @[RegFile.scala 65:20:@39249.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 65:20:@39249.4]
  wire  regs_426_io_enable; // @[RegFile.scala 65:20:@39249.4]
  wire  regs_427_clock; // @[RegFile.scala 65:20:@39263.4]
  wire  regs_427_reset; // @[RegFile.scala 65:20:@39263.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 65:20:@39263.4]
  wire  regs_427_io_reset; // @[RegFile.scala 65:20:@39263.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 65:20:@39263.4]
  wire  regs_427_io_enable; // @[RegFile.scala 65:20:@39263.4]
  wire  regs_428_clock; // @[RegFile.scala 65:20:@39277.4]
  wire  regs_428_reset; // @[RegFile.scala 65:20:@39277.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 65:20:@39277.4]
  wire  regs_428_io_reset; // @[RegFile.scala 65:20:@39277.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 65:20:@39277.4]
  wire  regs_428_io_enable; // @[RegFile.scala 65:20:@39277.4]
  wire  regs_429_clock; // @[RegFile.scala 65:20:@39291.4]
  wire  regs_429_reset; // @[RegFile.scala 65:20:@39291.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 65:20:@39291.4]
  wire  regs_429_io_reset; // @[RegFile.scala 65:20:@39291.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 65:20:@39291.4]
  wire  regs_429_io_enable; // @[RegFile.scala 65:20:@39291.4]
  wire  regs_430_clock; // @[RegFile.scala 65:20:@39305.4]
  wire  regs_430_reset; // @[RegFile.scala 65:20:@39305.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 65:20:@39305.4]
  wire  regs_430_io_reset; // @[RegFile.scala 65:20:@39305.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 65:20:@39305.4]
  wire  regs_430_io_enable; // @[RegFile.scala 65:20:@39305.4]
  wire  regs_431_clock; // @[RegFile.scala 65:20:@39319.4]
  wire  regs_431_reset; // @[RegFile.scala 65:20:@39319.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 65:20:@39319.4]
  wire  regs_431_io_reset; // @[RegFile.scala 65:20:@39319.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 65:20:@39319.4]
  wire  regs_431_io_enable; // @[RegFile.scala 65:20:@39319.4]
  wire  regs_432_clock; // @[RegFile.scala 65:20:@39333.4]
  wire  regs_432_reset; // @[RegFile.scala 65:20:@39333.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 65:20:@39333.4]
  wire  regs_432_io_reset; // @[RegFile.scala 65:20:@39333.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 65:20:@39333.4]
  wire  regs_432_io_enable; // @[RegFile.scala 65:20:@39333.4]
  wire  regs_433_clock; // @[RegFile.scala 65:20:@39347.4]
  wire  regs_433_reset; // @[RegFile.scala 65:20:@39347.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 65:20:@39347.4]
  wire  regs_433_io_reset; // @[RegFile.scala 65:20:@39347.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 65:20:@39347.4]
  wire  regs_433_io_enable; // @[RegFile.scala 65:20:@39347.4]
  wire  regs_434_clock; // @[RegFile.scala 65:20:@39361.4]
  wire  regs_434_reset; // @[RegFile.scala 65:20:@39361.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 65:20:@39361.4]
  wire  regs_434_io_reset; // @[RegFile.scala 65:20:@39361.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 65:20:@39361.4]
  wire  regs_434_io_enable; // @[RegFile.scala 65:20:@39361.4]
  wire  regs_435_clock; // @[RegFile.scala 65:20:@39375.4]
  wire  regs_435_reset; // @[RegFile.scala 65:20:@39375.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 65:20:@39375.4]
  wire  regs_435_io_reset; // @[RegFile.scala 65:20:@39375.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 65:20:@39375.4]
  wire  regs_435_io_enable; // @[RegFile.scala 65:20:@39375.4]
  wire  regs_436_clock; // @[RegFile.scala 65:20:@39389.4]
  wire  regs_436_reset; // @[RegFile.scala 65:20:@39389.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 65:20:@39389.4]
  wire  regs_436_io_reset; // @[RegFile.scala 65:20:@39389.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 65:20:@39389.4]
  wire  regs_436_io_enable; // @[RegFile.scala 65:20:@39389.4]
  wire  regs_437_clock; // @[RegFile.scala 65:20:@39403.4]
  wire  regs_437_reset; // @[RegFile.scala 65:20:@39403.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 65:20:@39403.4]
  wire  regs_437_io_reset; // @[RegFile.scala 65:20:@39403.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 65:20:@39403.4]
  wire  regs_437_io_enable; // @[RegFile.scala 65:20:@39403.4]
  wire  regs_438_clock; // @[RegFile.scala 65:20:@39417.4]
  wire  regs_438_reset; // @[RegFile.scala 65:20:@39417.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 65:20:@39417.4]
  wire  regs_438_io_reset; // @[RegFile.scala 65:20:@39417.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 65:20:@39417.4]
  wire  regs_438_io_enable; // @[RegFile.scala 65:20:@39417.4]
  wire  regs_439_clock; // @[RegFile.scala 65:20:@39431.4]
  wire  regs_439_reset; // @[RegFile.scala 65:20:@39431.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 65:20:@39431.4]
  wire  regs_439_io_reset; // @[RegFile.scala 65:20:@39431.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 65:20:@39431.4]
  wire  regs_439_io_enable; // @[RegFile.scala 65:20:@39431.4]
  wire  regs_440_clock; // @[RegFile.scala 65:20:@39445.4]
  wire  regs_440_reset; // @[RegFile.scala 65:20:@39445.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 65:20:@39445.4]
  wire  regs_440_io_reset; // @[RegFile.scala 65:20:@39445.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 65:20:@39445.4]
  wire  regs_440_io_enable; // @[RegFile.scala 65:20:@39445.4]
  wire  regs_441_clock; // @[RegFile.scala 65:20:@39459.4]
  wire  regs_441_reset; // @[RegFile.scala 65:20:@39459.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 65:20:@39459.4]
  wire  regs_441_io_reset; // @[RegFile.scala 65:20:@39459.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 65:20:@39459.4]
  wire  regs_441_io_enable; // @[RegFile.scala 65:20:@39459.4]
  wire  regs_442_clock; // @[RegFile.scala 65:20:@39473.4]
  wire  regs_442_reset; // @[RegFile.scala 65:20:@39473.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 65:20:@39473.4]
  wire  regs_442_io_reset; // @[RegFile.scala 65:20:@39473.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 65:20:@39473.4]
  wire  regs_442_io_enable; // @[RegFile.scala 65:20:@39473.4]
  wire  regs_443_clock; // @[RegFile.scala 65:20:@39487.4]
  wire  regs_443_reset; // @[RegFile.scala 65:20:@39487.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 65:20:@39487.4]
  wire  regs_443_io_reset; // @[RegFile.scala 65:20:@39487.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 65:20:@39487.4]
  wire  regs_443_io_enable; // @[RegFile.scala 65:20:@39487.4]
  wire  regs_444_clock; // @[RegFile.scala 65:20:@39501.4]
  wire  regs_444_reset; // @[RegFile.scala 65:20:@39501.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 65:20:@39501.4]
  wire  regs_444_io_reset; // @[RegFile.scala 65:20:@39501.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 65:20:@39501.4]
  wire  regs_444_io_enable; // @[RegFile.scala 65:20:@39501.4]
  wire  regs_445_clock; // @[RegFile.scala 65:20:@39515.4]
  wire  regs_445_reset; // @[RegFile.scala 65:20:@39515.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 65:20:@39515.4]
  wire  regs_445_io_reset; // @[RegFile.scala 65:20:@39515.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 65:20:@39515.4]
  wire  regs_445_io_enable; // @[RegFile.scala 65:20:@39515.4]
  wire  regs_446_clock; // @[RegFile.scala 65:20:@39529.4]
  wire  regs_446_reset; // @[RegFile.scala 65:20:@39529.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 65:20:@39529.4]
  wire  regs_446_io_reset; // @[RegFile.scala 65:20:@39529.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 65:20:@39529.4]
  wire  regs_446_io_enable; // @[RegFile.scala 65:20:@39529.4]
  wire  regs_447_clock; // @[RegFile.scala 65:20:@39543.4]
  wire  regs_447_reset; // @[RegFile.scala 65:20:@39543.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 65:20:@39543.4]
  wire  regs_447_io_reset; // @[RegFile.scala 65:20:@39543.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 65:20:@39543.4]
  wire  regs_447_io_enable; // @[RegFile.scala 65:20:@39543.4]
  wire  regs_448_clock; // @[RegFile.scala 65:20:@39557.4]
  wire  regs_448_reset; // @[RegFile.scala 65:20:@39557.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 65:20:@39557.4]
  wire  regs_448_io_reset; // @[RegFile.scala 65:20:@39557.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 65:20:@39557.4]
  wire  regs_448_io_enable; // @[RegFile.scala 65:20:@39557.4]
  wire  regs_449_clock; // @[RegFile.scala 65:20:@39571.4]
  wire  regs_449_reset; // @[RegFile.scala 65:20:@39571.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 65:20:@39571.4]
  wire  regs_449_io_reset; // @[RegFile.scala 65:20:@39571.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 65:20:@39571.4]
  wire  regs_449_io_enable; // @[RegFile.scala 65:20:@39571.4]
  wire  regs_450_clock; // @[RegFile.scala 65:20:@39585.4]
  wire  regs_450_reset; // @[RegFile.scala 65:20:@39585.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 65:20:@39585.4]
  wire  regs_450_io_reset; // @[RegFile.scala 65:20:@39585.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 65:20:@39585.4]
  wire  regs_450_io_enable; // @[RegFile.scala 65:20:@39585.4]
  wire  regs_451_clock; // @[RegFile.scala 65:20:@39599.4]
  wire  regs_451_reset; // @[RegFile.scala 65:20:@39599.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 65:20:@39599.4]
  wire  regs_451_io_reset; // @[RegFile.scala 65:20:@39599.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 65:20:@39599.4]
  wire  regs_451_io_enable; // @[RegFile.scala 65:20:@39599.4]
  wire  regs_452_clock; // @[RegFile.scala 65:20:@39613.4]
  wire  regs_452_reset; // @[RegFile.scala 65:20:@39613.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 65:20:@39613.4]
  wire  regs_452_io_reset; // @[RegFile.scala 65:20:@39613.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 65:20:@39613.4]
  wire  regs_452_io_enable; // @[RegFile.scala 65:20:@39613.4]
  wire  regs_453_clock; // @[RegFile.scala 65:20:@39627.4]
  wire  regs_453_reset; // @[RegFile.scala 65:20:@39627.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 65:20:@39627.4]
  wire  regs_453_io_reset; // @[RegFile.scala 65:20:@39627.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 65:20:@39627.4]
  wire  regs_453_io_enable; // @[RegFile.scala 65:20:@39627.4]
  wire  regs_454_clock; // @[RegFile.scala 65:20:@39641.4]
  wire  regs_454_reset; // @[RegFile.scala 65:20:@39641.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 65:20:@39641.4]
  wire  regs_454_io_reset; // @[RegFile.scala 65:20:@39641.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 65:20:@39641.4]
  wire  regs_454_io_enable; // @[RegFile.scala 65:20:@39641.4]
  wire  regs_455_clock; // @[RegFile.scala 65:20:@39655.4]
  wire  regs_455_reset; // @[RegFile.scala 65:20:@39655.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 65:20:@39655.4]
  wire  regs_455_io_reset; // @[RegFile.scala 65:20:@39655.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 65:20:@39655.4]
  wire  regs_455_io_enable; // @[RegFile.scala 65:20:@39655.4]
  wire  regs_456_clock; // @[RegFile.scala 65:20:@39669.4]
  wire  regs_456_reset; // @[RegFile.scala 65:20:@39669.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 65:20:@39669.4]
  wire  regs_456_io_reset; // @[RegFile.scala 65:20:@39669.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 65:20:@39669.4]
  wire  regs_456_io_enable; // @[RegFile.scala 65:20:@39669.4]
  wire  regs_457_clock; // @[RegFile.scala 65:20:@39683.4]
  wire  regs_457_reset; // @[RegFile.scala 65:20:@39683.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 65:20:@39683.4]
  wire  regs_457_io_reset; // @[RegFile.scala 65:20:@39683.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 65:20:@39683.4]
  wire  regs_457_io_enable; // @[RegFile.scala 65:20:@39683.4]
  wire  regs_458_clock; // @[RegFile.scala 65:20:@39697.4]
  wire  regs_458_reset; // @[RegFile.scala 65:20:@39697.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 65:20:@39697.4]
  wire  regs_458_io_reset; // @[RegFile.scala 65:20:@39697.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 65:20:@39697.4]
  wire  regs_458_io_enable; // @[RegFile.scala 65:20:@39697.4]
  wire  regs_459_clock; // @[RegFile.scala 65:20:@39711.4]
  wire  regs_459_reset; // @[RegFile.scala 65:20:@39711.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 65:20:@39711.4]
  wire  regs_459_io_reset; // @[RegFile.scala 65:20:@39711.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 65:20:@39711.4]
  wire  regs_459_io_enable; // @[RegFile.scala 65:20:@39711.4]
  wire  regs_460_clock; // @[RegFile.scala 65:20:@39725.4]
  wire  regs_460_reset; // @[RegFile.scala 65:20:@39725.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 65:20:@39725.4]
  wire  regs_460_io_reset; // @[RegFile.scala 65:20:@39725.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 65:20:@39725.4]
  wire  regs_460_io_enable; // @[RegFile.scala 65:20:@39725.4]
  wire  regs_461_clock; // @[RegFile.scala 65:20:@39739.4]
  wire  regs_461_reset; // @[RegFile.scala 65:20:@39739.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 65:20:@39739.4]
  wire  regs_461_io_reset; // @[RegFile.scala 65:20:@39739.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 65:20:@39739.4]
  wire  regs_461_io_enable; // @[RegFile.scala 65:20:@39739.4]
  wire  regs_462_clock; // @[RegFile.scala 65:20:@39753.4]
  wire  regs_462_reset; // @[RegFile.scala 65:20:@39753.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 65:20:@39753.4]
  wire  regs_462_io_reset; // @[RegFile.scala 65:20:@39753.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 65:20:@39753.4]
  wire  regs_462_io_enable; // @[RegFile.scala 65:20:@39753.4]
  wire  regs_463_clock; // @[RegFile.scala 65:20:@39767.4]
  wire  regs_463_reset; // @[RegFile.scala 65:20:@39767.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 65:20:@39767.4]
  wire  regs_463_io_reset; // @[RegFile.scala 65:20:@39767.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 65:20:@39767.4]
  wire  regs_463_io_enable; // @[RegFile.scala 65:20:@39767.4]
  wire  regs_464_clock; // @[RegFile.scala 65:20:@39781.4]
  wire  regs_464_reset; // @[RegFile.scala 65:20:@39781.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 65:20:@39781.4]
  wire  regs_464_io_reset; // @[RegFile.scala 65:20:@39781.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 65:20:@39781.4]
  wire  regs_464_io_enable; // @[RegFile.scala 65:20:@39781.4]
  wire  regs_465_clock; // @[RegFile.scala 65:20:@39795.4]
  wire  regs_465_reset; // @[RegFile.scala 65:20:@39795.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 65:20:@39795.4]
  wire  regs_465_io_reset; // @[RegFile.scala 65:20:@39795.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 65:20:@39795.4]
  wire  regs_465_io_enable; // @[RegFile.scala 65:20:@39795.4]
  wire  regs_466_clock; // @[RegFile.scala 65:20:@39809.4]
  wire  regs_466_reset; // @[RegFile.scala 65:20:@39809.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 65:20:@39809.4]
  wire  regs_466_io_reset; // @[RegFile.scala 65:20:@39809.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 65:20:@39809.4]
  wire  regs_466_io_enable; // @[RegFile.scala 65:20:@39809.4]
  wire  regs_467_clock; // @[RegFile.scala 65:20:@39823.4]
  wire  regs_467_reset; // @[RegFile.scala 65:20:@39823.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 65:20:@39823.4]
  wire  regs_467_io_reset; // @[RegFile.scala 65:20:@39823.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 65:20:@39823.4]
  wire  regs_467_io_enable; // @[RegFile.scala 65:20:@39823.4]
  wire  regs_468_clock; // @[RegFile.scala 65:20:@39837.4]
  wire  regs_468_reset; // @[RegFile.scala 65:20:@39837.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 65:20:@39837.4]
  wire  regs_468_io_reset; // @[RegFile.scala 65:20:@39837.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 65:20:@39837.4]
  wire  regs_468_io_enable; // @[RegFile.scala 65:20:@39837.4]
  wire  regs_469_clock; // @[RegFile.scala 65:20:@39851.4]
  wire  regs_469_reset; // @[RegFile.scala 65:20:@39851.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 65:20:@39851.4]
  wire  regs_469_io_reset; // @[RegFile.scala 65:20:@39851.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 65:20:@39851.4]
  wire  regs_469_io_enable; // @[RegFile.scala 65:20:@39851.4]
  wire  regs_470_clock; // @[RegFile.scala 65:20:@39865.4]
  wire  regs_470_reset; // @[RegFile.scala 65:20:@39865.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 65:20:@39865.4]
  wire  regs_470_io_reset; // @[RegFile.scala 65:20:@39865.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 65:20:@39865.4]
  wire  regs_470_io_enable; // @[RegFile.scala 65:20:@39865.4]
  wire  regs_471_clock; // @[RegFile.scala 65:20:@39879.4]
  wire  regs_471_reset; // @[RegFile.scala 65:20:@39879.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 65:20:@39879.4]
  wire  regs_471_io_reset; // @[RegFile.scala 65:20:@39879.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 65:20:@39879.4]
  wire  regs_471_io_enable; // @[RegFile.scala 65:20:@39879.4]
  wire  regs_472_clock; // @[RegFile.scala 65:20:@39893.4]
  wire  regs_472_reset; // @[RegFile.scala 65:20:@39893.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 65:20:@39893.4]
  wire  regs_472_io_reset; // @[RegFile.scala 65:20:@39893.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 65:20:@39893.4]
  wire  regs_472_io_enable; // @[RegFile.scala 65:20:@39893.4]
  wire  regs_473_clock; // @[RegFile.scala 65:20:@39907.4]
  wire  regs_473_reset; // @[RegFile.scala 65:20:@39907.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 65:20:@39907.4]
  wire  regs_473_io_reset; // @[RegFile.scala 65:20:@39907.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 65:20:@39907.4]
  wire  regs_473_io_enable; // @[RegFile.scala 65:20:@39907.4]
  wire  regs_474_clock; // @[RegFile.scala 65:20:@39921.4]
  wire  regs_474_reset; // @[RegFile.scala 65:20:@39921.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 65:20:@39921.4]
  wire  regs_474_io_reset; // @[RegFile.scala 65:20:@39921.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 65:20:@39921.4]
  wire  regs_474_io_enable; // @[RegFile.scala 65:20:@39921.4]
  wire  regs_475_clock; // @[RegFile.scala 65:20:@39935.4]
  wire  regs_475_reset; // @[RegFile.scala 65:20:@39935.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 65:20:@39935.4]
  wire  regs_475_io_reset; // @[RegFile.scala 65:20:@39935.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 65:20:@39935.4]
  wire  regs_475_io_enable; // @[RegFile.scala 65:20:@39935.4]
  wire  regs_476_clock; // @[RegFile.scala 65:20:@39949.4]
  wire  regs_476_reset; // @[RegFile.scala 65:20:@39949.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 65:20:@39949.4]
  wire  regs_476_io_reset; // @[RegFile.scala 65:20:@39949.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 65:20:@39949.4]
  wire  regs_476_io_enable; // @[RegFile.scala 65:20:@39949.4]
  wire  regs_477_clock; // @[RegFile.scala 65:20:@39963.4]
  wire  regs_477_reset; // @[RegFile.scala 65:20:@39963.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 65:20:@39963.4]
  wire  regs_477_io_reset; // @[RegFile.scala 65:20:@39963.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 65:20:@39963.4]
  wire  regs_477_io_enable; // @[RegFile.scala 65:20:@39963.4]
  wire  regs_478_clock; // @[RegFile.scala 65:20:@39977.4]
  wire  regs_478_reset; // @[RegFile.scala 65:20:@39977.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 65:20:@39977.4]
  wire  regs_478_io_reset; // @[RegFile.scala 65:20:@39977.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 65:20:@39977.4]
  wire  regs_478_io_enable; // @[RegFile.scala 65:20:@39977.4]
  wire  regs_479_clock; // @[RegFile.scala 65:20:@39991.4]
  wire  regs_479_reset; // @[RegFile.scala 65:20:@39991.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 65:20:@39991.4]
  wire  regs_479_io_reset; // @[RegFile.scala 65:20:@39991.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 65:20:@39991.4]
  wire  regs_479_io_enable; // @[RegFile.scala 65:20:@39991.4]
  wire  regs_480_clock; // @[RegFile.scala 65:20:@40005.4]
  wire  regs_480_reset; // @[RegFile.scala 65:20:@40005.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 65:20:@40005.4]
  wire  regs_480_io_reset; // @[RegFile.scala 65:20:@40005.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 65:20:@40005.4]
  wire  regs_480_io_enable; // @[RegFile.scala 65:20:@40005.4]
  wire  regs_481_clock; // @[RegFile.scala 65:20:@40019.4]
  wire  regs_481_reset; // @[RegFile.scala 65:20:@40019.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 65:20:@40019.4]
  wire  regs_481_io_reset; // @[RegFile.scala 65:20:@40019.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 65:20:@40019.4]
  wire  regs_481_io_enable; // @[RegFile.scala 65:20:@40019.4]
  wire  regs_482_clock; // @[RegFile.scala 65:20:@40033.4]
  wire  regs_482_reset; // @[RegFile.scala 65:20:@40033.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 65:20:@40033.4]
  wire  regs_482_io_reset; // @[RegFile.scala 65:20:@40033.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 65:20:@40033.4]
  wire  regs_482_io_enable; // @[RegFile.scala 65:20:@40033.4]
  wire  regs_483_clock; // @[RegFile.scala 65:20:@40047.4]
  wire  regs_483_reset; // @[RegFile.scala 65:20:@40047.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 65:20:@40047.4]
  wire  regs_483_io_reset; // @[RegFile.scala 65:20:@40047.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 65:20:@40047.4]
  wire  regs_483_io_enable; // @[RegFile.scala 65:20:@40047.4]
  wire  regs_484_clock; // @[RegFile.scala 65:20:@40061.4]
  wire  regs_484_reset; // @[RegFile.scala 65:20:@40061.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 65:20:@40061.4]
  wire  regs_484_io_reset; // @[RegFile.scala 65:20:@40061.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 65:20:@40061.4]
  wire  regs_484_io_enable; // @[RegFile.scala 65:20:@40061.4]
  wire  regs_485_clock; // @[RegFile.scala 65:20:@40075.4]
  wire  regs_485_reset; // @[RegFile.scala 65:20:@40075.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 65:20:@40075.4]
  wire  regs_485_io_reset; // @[RegFile.scala 65:20:@40075.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 65:20:@40075.4]
  wire  regs_485_io_enable; // @[RegFile.scala 65:20:@40075.4]
  wire  regs_486_clock; // @[RegFile.scala 65:20:@40089.4]
  wire  regs_486_reset; // @[RegFile.scala 65:20:@40089.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 65:20:@40089.4]
  wire  regs_486_io_reset; // @[RegFile.scala 65:20:@40089.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 65:20:@40089.4]
  wire  regs_486_io_enable; // @[RegFile.scala 65:20:@40089.4]
  wire  regs_487_clock; // @[RegFile.scala 65:20:@40103.4]
  wire  regs_487_reset; // @[RegFile.scala 65:20:@40103.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 65:20:@40103.4]
  wire  regs_487_io_reset; // @[RegFile.scala 65:20:@40103.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 65:20:@40103.4]
  wire  regs_487_io_enable; // @[RegFile.scala 65:20:@40103.4]
  wire  regs_488_clock; // @[RegFile.scala 65:20:@40117.4]
  wire  regs_488_reset; // @[RegFile.scala 65:20:@40117.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 65:20:@40117.4]
  wire  regs_488_io_reset; // @[RegFile.scala 65:20:@40117.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 65:20:@40117.4]
  wire  regs_488_io_enable; // @[RegFile.scala 65:20:@40117.4]
  wire  regs_489_clock; // @[RegFile.scala 65:20:@40131.4]
  wire  regs_489_reset; // @[RegFile.scala 65:20:@40131.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 65:20:@40131.4]
  wire  regs_489_io_reset; // @[RegFile.scala 65:20:@40131.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 65:20:@40131.4]
  wire  regs_489_io_enable; // @[RegFile.scala 65:20:@40131.4]
  wire  regs_490_clock; // @[RegFile.scala 65:20:@40145.4]
  wire  regs_490_reset; // @[RegFile.scala 65:20:@40145.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 65:20:@40145.4]
  wire  regs_490_io_reset; // @[RegFile.scala 65:20:@40145.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 65:20:@40145.4]
  wire  regs_490_io_enable; // @[RegFile.scala 65:20:@40145.4]
  wire  regs_491_clock; // @[RegFile.scala 65:20:@40159.4]
  wire  regs_491_reset; // @[RegFile.scala 65:20:@40159.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 65:20:@40159.4]
  wire  regs_491_io_reset; // @[RegFile.scala 65:20:@40159.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 65:20:@40159.4]
  wire  regs_491_io_enable; // @[RegFile.scala 65:20:@40159.4]
  wire  regs_492_clock; // @[RegFile.scala 65:20:@40173.4]
  wire  regs_492_reset; // @[RegFile.scala 65:20:@40173.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 65:20:@40173.4]
  wire  regs_492_io_reset; // @[RegFile.scala 65:20:@40173.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 65:20:@40173.4]
  wire  regs_492_io_enable; // @[RegFile.scala 65:20:@40173.4]
  wire  regs_493_clock; // @[RegFile.scala 65:20:@40187.4]
  wire  regs_493_reset; // @[RegFile.scala 65:20:@40187.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 65:20:@40187.4]
  wire  regs_493_io_reset; // @[RegFile.scala 65:20:@40187.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 65:20:@40187.4]
  wire  regs_493_io_enable; // @[RegFile.scala 65:20:@40187.4]
  wire  regs_494_clock; // @[RegFile.scala 65:20:@40201.4]
  wire  regs_494_reset; // @[RegFile.scala 65:20:@40201.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 65:20:@40201.4]
  wire  regs_494_io_reset; // @[RegFile.scala 65:20:@40201.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 65:20:@40201.4]
  wire  regs_494_io_enable; // @[RegFile.scala 65:20:@40201.4]
  wire  regs_495_clock; // @[RegFile.scala 65:20:@40215.4]
  wire  regs_495_reset; // @[RegFile.scala 65:20:@40215.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 65:20:@40215.4]
  wire  regs_495_io_reset; // @[RegFile.scala 65:20:@40215.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 65:20:@40215.4]
  wire  regs_495_io_enable; // @[RegFile.scala 65:20:@40215.4]
  wire  regs_496_clock; // @[RegFile.scala 65:20:@40229.4]
  wire  regs_496_reset; // @[RegFile.scala 65:20:@40229.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 65:20:@40229.4]
  wire  regs_496_io_reset; // @[RegFile.scala 65:20:@40229.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 65:20:@40229.4]
  wire  regs_496_io_enable; // @[RegFile.scala 65:20:@40229.4]
  wire  regs_497_clock; // @[RegFile.scala 65:20:@40243.4]
  wire  regs_497_reset; // @[RegFile.scala 65:20:@40243.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 65:20:@40243.4]
  wire  regs_497_io_reset; // @[RegFile.scala 65:20:@40243.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 65:20:@40243.4]
  wire  regs_497_io_enable; // @[RegFile.scala 65:20:@40243.4]
  wire  regs_498_clock; // @[RegFile.scala 65:20:@40257.4]
  wire  regs_498_reset; // @[RegFile.scala 65:20:@40257.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 65:20:@40257.4]
  wire  regs_498_io_reset; // @[RegFile.scala 65:20:@40257.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 65:20:@40257.4]
  wire  regs_498_io_enable; // @[RegFile.scala 65:20:@40257.4]
  wire  regs_499_clock; // @[RegFile.scala 65:20:@40271.4]
  wire  regs_499_reset; // @[RegFile.scala 65:20:@40271.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 65:20:@40271.4]
  wire  regs_499_io_reset; // @[RegFile.scala 65:20:@40271.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 65:20:@40271.4]
  wire  regs_499_io_enable; // @[RegFile.scala 65:20:@40271.4]
  wire  regs_500_clock; // @[RegFile.scala 65:20:@40285.4]
  wire  regs_500_reset; // @[RegFile.scala 65:20:@40285.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 65:20:@40285.4]
  wire  regs_500_io_reset; // @[RegFile.scala 65:20:@40285.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 65:20:@40285.4]
  wire  regs_500_io_enable; // @[RegFile.scala 65:20:@40285.4]
  wire  regs_501_clock; // @[RegFile.scala 65:20:@40299.4]
  wire  regs_501_reset; // @[RegFile.scala 65:20:@40299.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 65:20:@40299.4]
  wire  regs_501_io_reset; // @[RegFile.scala 65:20:@40299.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 65:20:@40299.4]
  wire  regs_501_io_enable; // @[RegFile.scala 65:20:@40299.4]
  wire  regs_502_clock; // @[RegFile.scala 65:20:@40313.4]
  wire  regs_502_reset; // @[RegFile.scala 65:20:@40313.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 65:20:@40313.4]
  wire  regs_502_io_reset; // @[RegFile.scala 65:20:@40313.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 65:20:@40313.4]
  wire  regs_502_io_enable; // @[RegFile.scala 65:20:@40313.4]
  FringeFF regs_0 ( // @[RegFile.scala 65:20:@33284.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 65:20:@33296.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 65:20:@33315.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 65:20:@33327.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 65:20:@33341.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 65:20:@33355.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 65:20:@33369.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 65:20:@33383.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 65:20:@33397.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 65:20:@33411.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 65:20:@33425.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 65:20:@33439.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 65:20:@33453.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 65:20:@33467.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 65:20:@33481.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 65:20:@33495.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 65:20:@33509.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 65:20:@33523.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 65:20:@33537.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 65:20:@33551.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 65:20:@33565.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 65:20:@33579.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 65:20:@33593.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 65:20:@33607.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 65:20:@33621.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 65:20:@33635.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 65:20:@33649.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 65:20:@33663.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 65:20:@33677.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 65:20:@33691.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 65:20:@33705.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 65:20:@33719.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 65:20:@33733.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 65:20:@33747.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 65:20:@33761.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 65:20:@33775.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 65:20:@33789.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 65:20:@33803.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 65:20:@33817.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 65:20:@33831.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 65:20:@33845.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 65:20:@33859.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 65:20:@33873.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 65:20:@33887.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 65:20:@33901.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 65:20:@33915.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 65:20:@33929.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 65:20:@33943.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 65:20:@33957.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 65:20:@33971.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 65:20:@33985.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 65:20:@33999.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 65:20:@34013.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 65:20:@34027.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 65:20:@34041.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 65:20:@34055.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 65:20:@34069.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 65:20:@34083.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 65:20:@34097.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 65:20:@34111.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 65:20:@34125.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 65:20:@34139.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 65:20:@34153.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 65:20:@34167.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 65:20:@34181.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 65:20:@34195.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 65:20:@34209.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 65:20:@34223.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 65:20:@34237.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 65:20:@34251.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 65:20:@34265.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 65:20:@34279.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 65:20:@34293.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 65:20:@34307.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 65:20:@34321.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 65:20:@34335.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 65:20:@34349.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 65:20:@34363.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 65:20:@34377.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 65:20:@34391.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 65:20:@34405.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 65:20:@34419.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 65:20:@34433.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 65:20:@34447.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 65:20:@34461.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 65:20:@34475.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 65:20:@34489.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 65:20:@34503.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 65:20:@34517.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 65:20:@34531.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 65:20:@34545.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 65:20:@34559.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 65:20:@34573.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 65:20:@34587.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 65:20:@34601.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 65:20:@34615.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 65:20:@34629.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 65:20:@34643.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 65:20:@34657.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 65:20:@34671.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 65:20:@34685.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 65:20:@34699.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 65:20:@34713.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 65:20:@34727.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 65:20:@34741.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 65:20:@34755.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 65:20:@34769.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 65:20:@34783.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 65:20:@34797.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 65:20:@34811.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 65:20:@34825.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 65:20:@34839.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 65:20:@34853.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 65:20:@34867.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 65:20:@34881.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 65:20:@34895.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 65:20:@34909.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 65:20:@34923.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 65:20:@34937.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 65:20:@34951.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 65:20:@34965.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 65:20:@34979.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 65:20:@34993.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 65:20:@35007.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 65:20:@35021.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 65:20:@35035.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 65:20:@35049.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 65:20:@35063.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 65:20:@35077.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 65:20:@35091.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 65:20:@35105.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 65:20:@35119.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 65:20:@35133.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 65:20:@35147.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 65:20:@35161.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 65:20:@35175.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 65:20:@35189.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 65:20:@35203.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 65:20:@35217.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 65:20:@35231.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 65:20:@35245.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 65:20:@35259.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 65:20:@35273.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 65:20:@35287.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 65:20:@35301.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 65:20:@35315.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 65:20:@35329.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 65:20:@35343.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 65:20:@35357.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 65:20:@35371.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 65:20:@35385.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 65:20:@35399.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 65:20:@35413.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 65:20:@35427.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 65:20:@35441.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 65:20:@35455.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 65:20:@35469.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 65:20:@35483.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 65:20:@35497.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 65:20:@35511.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 65:20:@35525.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 65:20:@35539.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 65:20:@35553.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 65:20:@35567.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 65:20:@35581.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 65:20:@35595.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 65:20:@35609.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 65:20:@35623.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 65:20:@35637.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 65:20:@35651.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 65:20:@35665.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 65:20:@35679.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 65:20:@35693.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 65:20:@35707.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 65:20:@35721.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 65:20:@35735.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 65:20:@35749.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 65:20:@35763.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 65:20:@35777.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 65:20:@35791.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 65:20:@35805.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 65:20:@35819.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 65:20:@35833.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 65:20:@35847.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 65:20:@35861.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 65:20:@35875.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 65:20:@35889.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 65:20:@35903.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 65:20:@35917.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 65:20:@35931.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 65:20:@35945.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 65:20:@35959.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 65:20:@35973.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 65:20:@35987.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 65:20:@36001.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 65:20:@36015.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 65:20:@36029.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 65:20:@36043.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 65:20:@36057.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 65:20:@36071.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 65:20:@36085.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 65:20:@36099.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 65:20:@36113.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 65:20:@36127.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 65:20:@36141.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 65:20:@36155.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 65:20:@36169.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 65:20:@36183.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 65:20:@36197.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 65:20:@36211.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 65:20:@36225.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 65:20:@36239.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 65:20:@36253.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 65:20:@36267.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 65:20:@36281.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 65:20:@36295.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 65:20:@36309.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 65:20:@36323.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 65:20:@36337.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 65:20:@36351.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 65:20:@36365.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 65:20:@36379.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 65:20:@36393.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 65:20:@36407.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 65:20:@36421.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 65:20:@36435.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 65:20:@36449.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 65:20:@36463.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 65:20:@36477.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 65:20:@36491.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 65:20:@36505.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 65:20:@36519.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 65:20:@36533.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 65:20:@36547.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 65:20:@36561.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 65:20:@36575.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 65:20:@36589.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 65:20:@36603.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 65:20:@36617.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 65:20:@36631.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 65:20:@36645.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 65:20:@36659.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 65:20:@36673.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 65:20:@36687.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 65:20:@36701.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 65:20:@36715.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 65:20:@36729.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 65:20:@36743.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 65:20:@36757.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 65:20:@36771.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 65:20:@36785.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 65:20:@36799.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 65:20:@36813.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 65:20:@36827.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 65:20:@36841.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 65:20:@36855.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 65:20:@36869.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 65:20:@36883.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 65:20:@36897.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 65:20:@36911.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 65:20:@36925.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 65:20:@36939.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 65:20:@36953.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 65:20:@36967.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 65:20:@36981.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 65:20:@36995.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 65:20:@37009.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 65:20:@37023.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 65:20:@37037.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 65:20:@37051.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 65:20:@37065.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 65:20:@37079.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 65:20:@37093.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 65:20:@37107.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 65:20:@37121.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 65:20:@37135.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 65:20:@37149.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 65:20:@37163.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 65:20:@37177.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 65:20:@37191.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 65:20:@37205.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 65:20:@37219.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 65:20:@37233.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 65:20:@37247.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 65:20:@37261.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 65:20:@37275.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 65:20:@37289.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 65:20:@37303.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 65:20:@37317.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 65:20:@37331.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 65:20:@37345.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 65:20:@37359.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 65:20:@37373.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 65:20:@37387.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 65:20:@37401.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 65:20:@37415.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 65:20:@37429.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 65:20:@37443.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 65:20:@37457.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 65:20:@37471.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 65:20:@37485.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 65:20:@37499.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 65:20:@37513.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 65:20:@37527.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 65:20:@37541.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 65:20:@37555.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 65:20:@37569.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 65:20:@37583.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 65:20:@37597.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 65:20:@37611.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 65:20:@37625.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 65:20:@37639.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 65:20:@37653.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 65:20:@37667.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 65:20:@37681.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 65:20:@37695.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 65:20:@37709.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 65:20:@37723.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 65:20:@37737.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 65:20:@37751.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 65:20:@37765.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 65:20:@37779.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 65:20:@37793.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 65:20:@37807.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 65:20:@37821.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 65:20:@37835.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 65:20:@37849.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 65:20:@37863.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 65:20:@37877.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 65:20:@37891.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 65:20:@37905.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 65:20:@37919.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 65:20:@37933.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 65:20:@37947.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 65:20:@37961.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 65:20:@37975.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 65:20:@37989.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 65:20:@38003.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 65:20:@38017.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 65:20:@38031.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 65:20:@38045.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 65:20:@38059.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 65:20:@38073.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 65:20:@38087.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 65:20:@38101.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 65:20:@38115.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 65:20:@38129.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 65:20:@38143.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 65:20:@38157.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 65:20:@38171.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 65:20:@38185.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 65:20:@38199.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 65:20:@38213.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 65:20:@38227.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 65:20:@38241.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 65:20:@38255.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 65:20:@38269.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 65:20:@38283.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 65:20:@38297.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 65:20:@38311.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 65:20:@38325.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 65:20:@38339.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 65:20:@38353.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 65:20:@38367.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 65:20:@38381.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 65:20:@38395.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 65:20:@38409.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 65:20:@38423.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 65:20:@38437.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 65:20:@38451.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 65:20:@38465.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 65:20:@38479.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 65:20:@38493.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 65:20:@38507.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 65:20:@38521.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 65:20:@38535.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 65:20:@38549.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 65:20:@38563.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 65:20:@38577.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 65:20:@38591.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 65:20:@38605.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 65:20:@38619.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 65:20:@38633.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 65:20:@38647.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 65:20:@38661.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 65:20:@38675.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 65:20:@38689.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 65:20:@38703.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 65:20:@38717.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 65:20:@38731.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 65:20:@38745.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 65:20:@38759.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 65:20:@38773.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 65:20:@38787.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 65:20:@38801.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 65:20:@38815.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 65:20:@38829.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 65:20:@38843.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 65:20:@38857.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 65:20:@38871.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 65:20:@38885.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 65:20:@38899.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 65:20:@38913.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 65:20:@38927.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 65:20:@38941.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 65:20:@38955.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 65:20:@38969.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 65:20:@38983.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 65:20:@38997.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 65:20:@39011.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 65:20:@39025.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 65:20:@39039.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 65:20:@39053.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 65:20:@39067.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 65:20:@39081.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 65:20:@39095.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 65:20:@39109.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 65:20:@39123.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 65:20:@39137.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 65:20:@39151.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 65:20:@39165.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 65:20:@39179.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 65:20:@39193.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 65:20:@39207.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 65:20:@39221.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 65:20:@39235.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 65:20:@39249.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 65:20:@39263.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 65:20:@39277.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 65:20:@39291.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 65:20:@39305.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 65:20:@39319.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 65:20:@39333.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 65:20:@39347.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 65:20:@39361.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 65:20:@39375.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 65:20:@39389.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 65:20:@39403.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 65:20:@39417.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 65:20:@39431.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 65:20:@39445.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 65:20:@39459.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 65:20:@39473.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 65:20:@39487.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 65:20:@39501.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 65:20:@39515.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 65:20:@39529.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 65:20:@39543.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 65:20:@39557.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 65:20:@39571.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 65:20:@39585.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 65:20:@39599.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 65:20:@39613.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 65:20:@39627.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 65:20:@39641.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 65:20:@39655.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 65:20:@39669.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 65:20:@39683.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 65:20:@39697.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 65:20:@39711.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 65:20:@39725.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 65:20:@39739.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 65:20:@39753.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 65:20:@39767.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 65:20:@39781.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 65:20:@39795.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 65:20:@39809.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 65:20:@39823.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 65:20:@39837.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 65:20:@39851.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 65:20:@39865.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 65:20:@39879.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 65:20:@39893.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 65:20:@39907.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 65:20:@39921.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 65:20:@39935.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 65:20:@39949.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 65:20:@39963.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 65:20:@39977.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 65:20:@39991.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 65:20:@40005.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 65:20:@40019.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 65:20:@40033.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 65:20:@40047.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 65:20:@40061.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 65:20:@40075.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 65:20:@40089.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 65:20:@40103.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 65:20:@40117.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 65:20:@40131.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 65:20:@40145.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 65:20:@40159.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 65:20:@40173.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 65:20:@40187.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 65:20:@40201.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 65:20:@40215.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 65:20:@40229.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 65:20:@40243.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 65:20:@40257.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 65:20:@40271.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 65:20:@40285.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 65:20:@40299.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 65:20:@40313.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 110:13:@41343.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 110:13:@41344.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 110:13:@41345.4]
  assign regs_0_clock = clock; // @[:@33285.4]
  assign regs_0_reset = reset; // @[:@33286.4 RegFile.scala 81:16:@33292.4]
  assign regs_0_io_in = 64'h0; // @[RegFile.scala 80:16:@33290.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 82:19:@33294.4]
  assign regs_0_io_enable = 1'h0; // @[RegFile.scala 79:20:@33289.4]
  assign regs_1_clock = clock; // @[:@33297.4]
  assign regs_1_reset = reset; // @[:@33298.4 RegFile.scala 69:16:@33310.4]
  assign regs_1_io_in = io_argOuts_0_bits; // @[RegFile.scala 68:16:@33308.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 71:19:@33313.4]
  assign regs_1_io_enable = io_argOuts_0_valid; // @[RegFile.scala 67:20:@33304.4]
  assign regs_2_clock = clock; // @[:@33316.4]
  assign regs_2_reset = reset; // @[:@33317.4 RegFile.scala 81:16:@33323.4]
  assign regs_2_io_in = 64'h0; // @[RegFile.scala 80:16:@33321.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 82:19:@33325.4]
  assign regs_2_io_enable = 1'h0; // @[RegFile.scala 79:20:@33320.4]
  assign regs_3_clock = clock; // @[:@33328.4]
  assign regs_3_reset = io_reset; // @[:@33329.4 RegFile.scala 75:16:@33336.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : 64'h0; // @[RegFile.scala 74:16:@33335.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 77:19:@33339.4]
  assign regs_3_io_enable = io_argOuts_1_valid; // @[RegFile.scala 73:20:@33333.4]
  assign regs_4_clock = clock; // @[:@33342.4]
  assign regs_4_reset = io_reset; // @[:@33343.4 RegFile.scala 75:16:@33350.4]
  assign regs_4_io_in = 64'h0; // @[RegFile.scala 74:16:@33349.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 77:19:@33353.4]
  assign regs_4_io_enable = 1'h1; // @[RegFile.scala 73:20:@33347.4]
  assign regs_5_clock = clock; // @[:@33356.4]
  assign regs_5_reset = io_reset; // @[:@33357.4 RegFile.scala 75:16:@33364.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 74:16:@33363.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 77:19:@33367.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 73:20:@33361.4]
  assign regs_6_clock = clock; // @[:@33370.4]
  assign regs_6_reset = io_reset; // @[:@33371.4 RegFile.scala 75:16:@33378.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 74:16:@33377.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 77:19:@33381.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 73:20:@33375.4]
  assign regs_7_clock = clock; // @[:@33384.4]
  assign regs_7_reset = io_reset; // @[:@33385.4 RegFile.scala 75:16:@33392.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 74:16:@33391.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 77:19:@33395.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 73:20:@33389.4]
  assign regs_8_clock = clock; // @[:@33398.4]
  assign regs_8_reset = io_reset; // @[:@33399.4 RegFile.scala 75:16:@33406.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 74:16:@33405.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 77:19:@33409.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 73:20:@33403.4]
  assign regs_9_clock = clock; // @[:@33412.4]
  assign regs_9_reset = io_reset; // @[:@33413.4 RegFile.scala 75:16:@33420.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 74:16:@33419.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 77:19:@33423.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 73:20:@33417.4]
  assign regs_10_clock = clock; // @[:@33426.4]
  assign regs_10_reset = io_reset; // @[:@33427.4 RegFile.scala 75:16:@33434.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 74:16:@33433.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 77:19:@33437.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 73:20:@33431.4]
  assign regs_11_clock = clock; // @[:@33440.4]
  assign regs_11_reset = io_reset; // @[:@33441.4 RegFile.scala 75:16:@33448.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 74:16:@33447.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 77:19:@33451.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 73:20:@33445.4]
  assign regs_12_clock = clock; // @[:@33454.4]
  assign regs_12_reset = io_reset; // @[:@33455.4 RegFile.scala 75:16:@33462.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 74:16:@33461.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 77:19:@33465.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 73:20:@33459.4]
  assign regs_13_clock = clock; // @[:@33468.4]
  assign regs_13_reset = io_reset; // @[:@33469.4 RegFile.scala 75:16:@33476.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 74:16:@33475.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 77:19:@33479.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 73:20:@33473.4]
  assign regs_14_clock = clock; // @[:@33482.4]
  assign regs_14_reset = io_reset; // @[:@33483.4 RegFile.scala 75:16:@33490.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 74:16:@33489.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 77:19:@33493.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 73:20:@33487.4]
  assign regs_15_clock = clock; // @[:@33496.4]
  assign regs_15_reset = io_reset; // @[:@33497.4 RegFile.scala 75:16:@33504.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 74:16:@33503.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 77:19:@33507.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 73:20:@33501.4]
  assign regs_16_clock = clock; // @[:@33510.4]
  assign regs_16_reset = io_reset; // @[:@33511.4 RegFile.scala 75:16:@33518.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 74:16:@33517.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 77:19:@33521.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 73:20:@33515.4]
  assign regs_17_clock = clock; // @[:@33524.4]
  assign regs_17_reset = io_reset; // @[:@33525.4 RegFile.scala 75:16:@33532.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 74:16:@33531.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 77:19:@33535.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 73:20:@33529.4]
  assign regs_18_clock = clock; // @[:@33538.4]
  assign regs_18_reset = io_reset; // @[:@33539.4 RegFile.scala 75:16:@33546.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 74:16:@33545.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 77:19:@33549.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 73:20:@33543.4]
  assign regs_19_clock = clock; // @[:@33552.4]
  assign regs_19_reset = io_reset; // @[:@33553.4 RegFile.scala 75:16:@33560.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 74:16:@33559.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 77:19:@33563.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 73:20:@33557.4]
  assign regs_20_clock = clock; // @[:@33566.4]
  assign regs_20_reset = io_reset; // @[:@33567.4 RegFile.scala 75:16:@33574.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 74:16:@33573.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 77:19:@33577.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 73:20:@33571.4]
  assign regs_21_clock = clock; // @[:@33580.4]
  assign regs_21_reset = io_reset; // @[:@33581.4 RegFile.scala 75:16:@33588.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 74:16:@33587.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 77:19:@33591.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 73:20:@33585.4]
  assign regs_22_clock = clock; // @[:@33594.4]
  assign regs_22_reset = io_reset; // @[:@33595.4 RegFile.scala 75:16:@33602.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 74:16:@33601.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 77:19:@33605.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 73:20:@33599.4]
  assign regs_23_clock = clock; // @[:@33608.4]
  assign regs_23_reset = io_reset; // @[:@33609.4 RegFile.scala 75:16:@33616.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 74:16:@33615.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 77:19:@33619.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 73:20:@33613.4]
  assign regs_24_clock = clock; // @[:@33622.4]
  assign regs_24_reset = io_reset; // @[:@33623.4 RegFile.scala 75:16:@33630.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 74:16:@33629.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 77:19:@33633.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 73:20:@33627.4]
  assign regs_25_clock = clock; // @[:@33636.4]
  assign regs_25_reset = io_reset; // @[:@33637.4 RegFile.scala 75:16:@33644.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 74:16:@33643.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 77:19:@33647.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 73:20:@33641.4]
  assign regs_26_clock = clock; // @[:@33650.4]
  assign regs_26_reset = io_reset; // @[:@33651.4 RegFile.scala 75:16:@33658.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 74:16:@33657.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 77:19:@33661.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 73:20:@33655.4]
  assign regs_27_clock = clock; // @[:@33664.4]
  assign regs_27_reset = io_reset; // @[:@33665.4 RegFile.scala 75:16:@33672.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 74:16:@33671.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 77:19:@33675.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 73:20:@33669.4]
  assign regs_28_clock = clock; // @[:@33678.4]
  assign regs_28_reset = io_reset; // @[:@33679.4 RegFile.scala 75:16:@33686.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 74:16:@33685.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 77:19:@33689.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 73:20:@33683.4]
  assign regs_29_clock = clock; // @[:@33692.4]
  assign regs_29_reset = io_reset; // @[:@33693.4 RegFile.scala 75:16:@33700.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 74:16:@33699.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 77:19:@33703.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 73:20:@33697.4]
  assign regs_30_clock = clock; // @[:@33706.4]
  assign regs_30_reset = io_reset; // @[:@33707.4 RegFile.scala 75:16:@33714.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 74:16:@33713.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 77:19:@33717.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 73:20:@33711.4]
  assign regs_31_clock = clock; // @[:@33720.4]
  assign regs_31_reset = io_reset; // @[:@33721.4 RegFile.scala 75:16:@33728.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 74:16:@33727.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 77:19:@33731.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 73:20:@33725.4]
  assign regs_32_clock = clock; // @[:@33734.4]
  assign regs_32_reset = io_reset; // @[:@33735.4 RegFile.scala 75:16:@33742.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 74:16:@33741.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 77:19:@33745.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 73:20:@33739.4]
  assign regs_33_clock = clock; // @[:@33748.4]
  assign regs_33_reset = io_reset; // @[:@33749.4 RegFile.scala 75:16:@33756.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 74:16:@33755.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 77:19:@33759.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 73:20:@33753.4]
  assign regs_34_clock = clock; // @[:@33762.4]
  assign regs_34_reset = io_reset; // @[:@33763.4 RegFile.scala 75:16:@33770.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 74:16:@33769.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 77:19:@33773.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 73:20:@33767.4]
  assign regs_35_clock = clock; // @[:@33776.4]
  assign regs_35_reset = io_reset; // @[:@33777.4 RegFile.scala 75:16:@33784.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 74:16:@33783.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 77:19:@33787.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 73:20:@33781.4]
  assign regs_36_clock = clock; // @[:@33790.4]
  assign regs_36_reset = io_reset; // @[:@33791.4 RegFile.scala 75:16:@33798.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 74:16:@33797.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 77:19:@33801.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 73:20:@33795.4]
  assign regs_37_clock = clock; // @[:@33804.4]
  assign regs_37_reset = io_reset; // @[:@33805.4 RegFile.scala 75:16:@33812.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 74:16:@33811.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 77:19:@33815.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 73:20:@33809.4]
  assign regs_38_clock = clock; // @[:@33818.4]
  assign regs_38_reset = io_reset; // @[:@33819.4 RegFile.scala 75:16:@33826.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 74:16:@33825.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 77:19:@33829.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 73:20:@33823.4]
  assign regs_39_clock = clock; // @[:@33832.4]
  assign regs_39_reset = io_reset; // @[:@33833.4 RegFile.scala 75:16:@33840.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 74:16:@33839.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 77:19:@33843.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 73:20:@33837.4]
  assign regs_40_clock = clock; // @[:@33846.4]
  assign regs_40_reset = io_reset; // @[:@33847.4 RegFile.scala 75:16:@33854.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 74:16:@33853.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 77:19:@33857.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 73:20:@33851.4]
  assign regs_41_clock = clock; // @[:@33860.4]
  assign regs_41_reset = io_reset; // @[:@33861.4 RegFile.scala 75:16:@33868.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 74:16:@33867.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 77:19:@33871.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 73:20:@33865.4]
  assign regs_42_clock = clock; // @[:@33874.4]
  assign regs_42_reset = io_reset; // @[:@33875.4 RegFile.scala 75:16:@33882.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 74:16:@33881.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 77:19:@33885.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 73:20:@33879.4]
  assign regs_43_clock = clock; // @[:@33888.4]
  assign regs_43_reset = io_reset; // @[:@33889.4 RegFile.scala 75:16:@33896.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 74:16:@33895.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 77:19:@33899.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 73:20:@33893.4]
  assign regs_44_clock = clock; // @[:@33902.4]
  assign regs_44_reset = io_reset; // @[:@33903.4 RegFile.scala 75:16:@33910.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 74:16:@33909.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 77:19:@33913.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 73:20:@33907.4]
  assign regs_45_clock = clock; // @[:@33916.4]
  assign regs_45_reset = io_reset; // @[:@33917.4 RegFile.scala 75:16:@33924.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 74:16:@33923.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 77:19:@33927.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 73:20:@33921.4]
  assign regs_46_clock = clock; // @[:@33930.4]
  assign regs_46_reset = io_reset; // @[:@33931.4 RegFile.scala 75:16:@33938.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 74:16:@33937.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 77:19:@33941.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 73:20:@33935.4]
  assign regs_47_clock = clock; // @[:@33944.4]
  assign regs_47_reset = io_reset; // @[:@33945.4 RegFile.scala 75:16:@33952.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 74:16:@33951.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 77:19:@33955.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 73:20:@33949.4]
  assign regs_48_clock = clock; // @[:@33958.4]
  assign regs_48_reset = io_reset; // @[:@33959.4 RegFile.scala 75:16:@33966.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 74:16:@33965.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 77:19:@33969.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 73:20:@33963.4]
  assign regs_49_clock = clock; // @[:@33972.4]
  assign regs_49_reset = io_reset; // @[:@33973.4 RegFile.scala 75:16:@33980.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 74:16:@33979.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 77:19:@33983.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 73:20:@33977.4]
  assign regs_50_clock = clock; // @[:@33986.4]
  assign regs_50_reset = io_reset; // @[:@33987.4 RegFile.scala 75:16:@33994.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 74:16:@33993.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 77:19:@33997.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 73:20:@33991.4]
  assign regs_51_clock = clock; // @[:@34000.4]
  assign regs_51_reset = io_reset; // @[:@34001.4 RegFile.scala 75:16:@34008.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 74:16:@34007.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 77:19:@34011.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 73:20:@34005.4]
  assign regs_52_clock = clock; // @[:@34014.4]
  assign regs_52_reset = io_reset; // @[:@34015.4 RegFile.scala 75:16:@34022.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 74:16:@34021.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 77:19:@34025.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 73:20:@34019.4]
  assign regs_53_clock = clock; // @[:@34028.4]
  assign regs_53_reset = io_reset; // @[:@34029.4 RegFile.scala 75:16:@34036.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 74:16:@34035.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 77:19:@34039.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 73:20:@34033.4]
  assign regs_54_clock = clock; // @[:@34042.4]
  assign regs_54_reset = io_reset; // @[:@34043.4 RegFile.scala 75:16:@34050.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 74:16:@34049.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 77:19:@34053.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 73:20:@34047.4]
  assign regs_55_clock = clock; // @[:@34056.4]
  assign regs_55_reset = io_reset; // @[:@34057.4 RegFile.scala 75:16:@34064.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 74:16:@34063.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 77:19:@34067.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 73:20:@34061.4]
  assign regs_56_clock = clock; // @[:@34070.4]
  assign regs_56_reset = io_reset; // @[:@34071.4 RegFile.scala 75:16:@34078.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 74:16:@34077.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 77:19:@34081.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 73:20:@34075.4]
  assign regs_57_clock = clock; // @[:@34084.4]
  assign regs_57_reset = io_reset; // @[:@34085.4 RegFile.scala 75:16:@34092.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 74:16:@34091.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 77:19:@34095.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 73:20:@34089.4]
  assign regs_58_clock = clock; // @[:@34098.4]
  assign regs_58_reset = io_reset; // @[:@34099.4 RegFile.scala 75:16:@34106.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 74:16:@34105.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 77:19:@34109.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 73:20:@34103.4]
  assign regs_59_clock = clock; // @[:@34112.4]
  assign regs_59_reset = io_reset; // @[:@34113.4 RegFile.scala 75:16:@34120.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 74:16:@34119.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 77:19:@34123.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 73:20:@34117.4]
  assign regs_60_clock = clock; // @[:@34126.4]
  assign regs_60_reset = io_reset; // @[:@34127.4 RegFile.scala 75:16:@34134.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 74:16:@34133.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 77:19:@34137.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 73:20:@34131.4]
  assign regs_61_clock = clock; // @[:@34140.4]
  assign regs_61_reset = io_reset; // @[:@34141.4 RegFile.scala 75:16:@34148.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 74:16:@34147.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 77:19:@34151.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 73:20:@34145.4]
  assign regs_62_clock = clock; // @[:@34154.4]
  assign regs_62_reset = io_reset; // @[:@34155.4 RegFile.scala 75:16:@34162.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 74:16:@34161.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 77:19:@34165.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 73:20:@34159.4]
  assign regs_63_clock = clock; // @[:@34168.4]
  assign regs_63_reset = io_reset; // @[:@34169.4 RegFile.scala 75:16:@34176.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 74:16:@34175.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 77:19:@34179.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 73:20:@34173.4]
  assign regs_64_clock = clock; // @[:@34182.4]
  assign regs_64_reset = io_reset; // @[:@34183.4 RegFile.scala 75:16:@34190.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 74:16:@34189.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 77:19:@34193.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 73:20:@34187.4]
  assign regs_65_clock = clock; // @[:@34196.4]
  assign regs_65_reset = io_reset; // @[:@34197.4 RegFile.scala 75:16:@34204.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 74:16:@34203.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 77:19:@34207.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 73:20:@34201.4]
  assign regs_66_clock = clock; // @[:@34210.4]
  assign regs_66_reset = io_reset; // @[:@34211.4 RegFile.scala 75:16:@34218.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 74:16:@34217.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 77:19:@34221.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 73:20:@34215.4]
  assign regs_67_clock = clock; // @[:@34224.4]
  assign regs_67_reset = io_reset; // @[:@34225.4 RegFile.scala 75:16:@34232.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 74:16:@34231.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 77:19:@34235.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 73:20:@34229.4]
  assign regs_68_clock = clock; // @[:@34238.4]
  assign regs_68_reset = io_reset; // @[:@34239.4 RegFile.scala 75:16:@34246.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 74:16:@34245.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 77:19:@34249.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 73:20:@34243.4]
  assign regs_69_clock = clock; // @[:@34252.4]
  assign regs_69_reset = io_reset; // @[:@34253.4 RegFile.scala 75:16:@34260.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 74:16:@34259.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 77:19:@34263.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 73:20:@34257.4]
  assign regs_70_clock = clock; // @[:@34266.4]
  assign regs_70_reset = io_reset; // @[:@34267.4 RegFile.scala 75:16:@34274.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 74:16:@34273.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 77:19:@34277.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 73:20:@34271.4]
  assign regs_71_clock = clock; // @[:@34280.4]
  assign regs_71_reset = io_reset; // @[:@34281.4 RegFile.scala 75:16:@34288.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 74:16:@34287.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 77:19:@34291.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 73:20:@34285.4]
  assign regs_72_clock = clock; // @[:@34294.4]
  assign regs_72_reset = io_reset; // @[:@34295.4 RegFile.scala 75:16:@34302.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 74:16:@34301.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 77:19:@34305.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 73:20:@34299.4]
  assign regs_73_clock = clock; // @[:@34308.4]
  assign regs_73_reset = io_reset; // @[:@34309.4 RegFile.scala 75:16:@34316.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 74:16:@34315.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 77:19:@34319.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 73:20:@34313.4]
  assign regs_74_clock = clock; // @[:@34322.4]
  assign regs_74_reset = io_reset; // @[:@34323.4 RegFile.scala 75:16:@34330.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 74:16:@34329.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 77:19:@34333.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 73:20:@34327.4]
  assign regs_75_clock = clock; // @[:@34336.4]
  assign regs_75_reset = io_reset; // @[:@34337.4 RegFile.scala 75:16:@34344.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 74:16:@34343.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 77:19:@34347.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 73:20:@34341.4]
  assign regs_76_clock = clock; // @[:@34350.4]
  assign regs_76_reset = io_reset; // @[:@34351.4 RegFile.scala 75:16:@34358.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 74:16:@34357.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 77:19:@34361.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 73:20:@34355.4]
  assign regs_77_clock = clock; // @[:@34364.4]
  assign regs_77_reset = io_reset; // @[:@34365.4 RegFile.scala 75:16:@34372.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 74:16:@34371.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 77:19:@34375.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 73:20:@34369.4]
  assign regs_78_clock = clock; // @[:@34378.4]
  assign regs_78_reset = io_reset; // @[:@34379.4 RegFile.scala 75:16:@34386.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 74:16:@34385.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 77:19:@34389.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 73:20:@34383.4]
  assign regs_79_clock = clock; // @[:@34392.4]
  assign regs_79_reset = io_reset; // @[:@34393.4 RegFile.scala 75:16:@34400.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 74:16:@34399.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 77:19:@34403.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 73:20:@34397.4]
  assign regs_80_clock = clock; // @[:@34406.4]
  assign regs_80_reset = io_reset; // @[:@34407.4 RegFile.scala 75:16:@34414.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 74:16:@34413.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 77:19:@34417.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 73:20:@34411.4]
  assign regs_81_clock = clock; // @[:@34420.4]
  assign regs_81_reset = io_reset; // @[:@34421.4 RegFile.scala 75:16:@34428.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 74:16:@34427.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 77:19:@34431.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 73:20:@34425.4]
  assign regs_82_clock = clock; // @[:@34434.4]
  assign regs_82_reset = io_reset; // @[:@34435.4 RegFile.scala 75:16:@34442.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 74:16:@34441.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 77:19:@34445.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 73:20:@34439.4]
  assign regs_83_clock = clock; // @[:@34448.4]
  assign regs_83_reset = io_reset; // @[:@34449.4 RegFile.scala 75:16:@34456.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 74:16:@34455.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 77:19:@34459.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 73:20:@34453.4]
  assign regs_84_clock = clock; // @[:@34462.4]
  assign regs_84_reset = io_reset; // @[:@34463.4 RegFile.scala 75:16:@34470.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 74:16:@34469.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 77:19:@34473.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 73:20:@34467.4]
  assign regs_85_clock = clock; // @[:@34476.4]
  assign regs_85_reset = io_reset; // @[:@34477.4 RegFile.scala 75:16:@34484.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 74:16:@34483.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 77:19:@34487.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 73:20:@34481.4]
  assign regs_86_clock = clock; // @[:@34490.4]
  assign regs_86_reset = io_reset; // @[:@34491.4 RegFile.scala 75:16:@34498.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 74:16:@34497.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 77:19:@34501.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 73:20:@34495.4]
  assign regs_87_clock = clock; // @[:@34504.4]
  assign regs_87_reset = io_reset; // @[:@34505.4 RegFile.scala 75:16:@34512.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 74:16:@34511.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 77:19:@34515.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 73:20:@34509.4]
  assign regs_88_clock = clock; // @[:@34518.4]
  assign regs_88_reset = io_reset; // @[:@34519.4 RegFile.scala 75:16:@34526.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 74:16:@34525.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 77:19:@34529.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 73:20:@34523.4]
  assign regs_89_clock = clock; // @[:@34532.4]
  assign regs_89_reset = io_reset; // @[:@34533.4 RegFile.scala 75:16:@34540.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 74:16:@34539.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 77:19:@34543.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 73:20:@34537.4]
  assign regs_90_clock = clock; // @[:@34546.4]
  assign regs_90_reset = io_reset; // @[:@34547.4 RegFile.scala 75:16:@34554.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 74:16:@34553.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 77:19:@34557.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 73:20:@34551.4]
  assign regs_91_clock = clock; // @[:@34560.4]
  assign regs_91_reset = io_reset; // @[:@34561.4 RegFile.scala 75:16:@34568.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 74:16:@34567.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 77:19:@34571.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 73:20:@34565.4]
  assign regs_92_clock = clock; // @[:@34574.4]
  assign regs_92_reset = io_reset; // @[:@34575.4 RegFile.scala 75:16:@34582.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 74:16:@34581.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 77:19:@34585.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 73:20:@34579.4]
  assign regs_93_clock = clock; // @[:@34588.4]
  assign regs_93_reset = io_reset; // @[:@34589.4 RegFile.scala 75:16:@34596.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 74:16:@34595.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 77:19:@34599.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 73:20:@34593.4]
  assign regs_94_clock = clock; // @[:@34602.4]
  assign regs_94_reset = io_reset; // @[:@34603.4 RegFile.scala 75:16:@34610.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 74:16:@34609.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 77:19:@34613.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 73:20:@34607.4]
  assign regs_95_clock = clock; // @[:@34616.4]
  assign regs_95_reset = io_reset; // @[:@34617.4 RegFile.scala 75:16:@34624.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 74:16:@34623.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 77:19:@34627.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 73:20:@34621.4]
  assign regs_96_clock = clock; // @[:@34630.4]
  assign regs_96_reset = io_reset; // @[:@34631.4 RegFile.scala 75:16:@34638.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 74:16:@34637.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 77:19:@34641.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 73:20:@34635.4]
  assign regs_97_clock = clock; // @[:@34644.4]
  assign regs_97_reset = io_reset; // @[:@34645.4 RegFile.scala 75:16:@34652.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 74:16:@34651.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 77:19:@34655.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 73:20:@34649.4]
  assign regs_98_clock = clock; // @[:@34658.4]
  assign regs_98_reset = io_reset; // @[:@34659.4 RegFile.scala 75:16:@34666.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 74:16:@34665.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 77:19:@34669.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 73:20:@34663.4]
  assign regs_99_clock = clock; // @[:@34672.4]
  assign regs_99_reset = io_reset; // @[:@34673.4 RegFile.scala 75:16:@34680.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 74:16:@34679.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 77:19:@34683.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 73:20:@34677.4]
  assign regs_100_clock = clock; // @[:@34686.4]
  assign regs_100_reset = io_reset; // @[:@34687.4 RegFile.scala 75:16:@34694.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 74:16:@34693.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 77:19:@34697.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 73:20:@34691.4]
  assign regs_101_clock = clock; // @[:@34700.4]
  assign regs_101_reset = io_reset; // @[:@34701.4 RegFile.scala 75:16:@34708.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 74:16:@34707.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 77:19:@34711.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 73:20:@34705.4]
  assign regs_102_clock = clock; // @[:@34714.4]
  assign regs_102_reset = io_reset; // @[:@34715.4 RegFile.scala 75:16:@34722.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 74:16:@34721.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 77:19:@34725.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 73:20:@34719.4]
  assign regs_103_clock = clock; // @[:@34728.4]
  assign regs_103_reset = io_reset; // @[:@34729.4 RegFile.scala 75:16:@34736.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 74:16:@34735.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 77:19:@34739.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 73:20:@34733.4]
  assign regs_104_clock = clock; // @[:@34742.4]
  assign regs_104_reset = io_reset; // @[:@34743.4 RegFile.scala 75:16:@34750.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 74:16:@34749.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 77:19:@34753.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 73:20:@34747.4]
  assign regs_105_clock = clock; // @[:@34756.4]
  assign regs_105_reset = io_reset; // @[:@34757.4 RegFile.scala 75:16:@34764.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 74:16:@34763.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 77:19:@34767.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 73:20:@34761.4]
  assign regs_106_clock = clock; // @[:@34770.4]
  assign regs_106_reset = io_reset; // @[:@34771.4 RegFile.scala 75:16:@34778.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 74:16:@34777.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 77:19:@34781.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 73:20:@34775.4]
  assign regs_107_clock = clock; // @[:@34784.4]
  assign regs_107_reset = io_reset; // @[:@34785.4 RegFile.scala 75:16:@34792.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 74:16:@34791.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 77:19:@34795.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 73:20:@34789.4]
  assign regs_108_clock = clock; // @[:@34798.4]
  assign regs_108_reset = io_reset; // @[:@34799.4 RegFile.scala 75:16:@34806.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 74:16:@34805.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 77:19:@34809.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 73:20:@34803.4]
  assign regs_109_clock = clock; // @[:@34812.4]
  assign regs_109_reset = io_reset; // @[:@34813.4 RegFile.scala 75:16:@34820.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 74:16:@34819.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 77:19:@34823.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 73:20:@34817.4]
  assign regs_110_clock = clock; // @[:@34826.4]
  assign regs_110_reset = io_reset; // @[:@34827.4 RegFile.scala 75:16:@34834.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 74:16:@34833.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 77:19:@34837.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 73:20:@34831.4]
  assign regs_111_clock = clock; // @[:@34840.4]
  assign regs_111_reset = io_reset; // @[:@34841.4 RegFile.scala 75:16:@34848.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 74:16:@34847.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 77:19:@34851.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 73:20:@34845.4]
  assign regs_112_clock = clock; // @[:@34854.4]
  assign regs_112_reset = io_reset; // @[:@34855.4 RegFile.scala 75:16:@34862.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 74:16:@34861.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 77:19:@34865.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 73:20:@34859.4]
  assign regs_113_clock = clock; // @[:@34868.4]
  assign regs_113_reset = io_reset; // @[:@34869.4 RegFile.scala 75:16:@34876.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 74:16:@34875.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 77:19:@34879.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 73:20:@34873.4]
  assign regs_114_clock = clock; // @[:@34882.4]
  assign regs_114_reset = io_reset; // @[:@34883.4 RegFile.scala 75:16:@34890.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 74:16:@34889.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 77:19:@34893.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 73:20:@34887.4]
  assign regs_115_clock = clock; // @[:@34896.4]
  assign regs_115_reset = io_reset; // @[:@34897.4 RegFile.scala 75:16:@34904.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 74:16:@34903.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 77:19:@34907.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 73:20:@34901.4]
  assign regs_116_clock = clock; // @[:@34910.4]
  assign regs_116_reset = io_reset; // @[:@34911.4 RegFile.scala 75:16:@34918.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 74:16:@34917.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 77:19:@34921.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 73:20:@34915.4]
  assign regs_117_clock = clock; // @[:@34924.4]
  assign regs_117_reset = io_reset; // @[:@34925.4 RegFile.scala 75:16:@34932.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 74:16:@34931.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 77:19:@34935.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 73:20:@34929.4]
  assign regs_118_clock = clock; // @[:@34938.4]
  assign regs_118_reset = io_reset; // @[:@34939.4 RegFile.scala 75:16:@34946.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 74:16:@34945.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 77:19:@34949.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 73:20:@34943.4]
  assign regs_119_clock = clock; // @[:@34952.4]
  assign regs_119_reset = io_reset; // @[:@34953.4 RegFile.scala 75:16:@34960.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 74:16:@34959.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 77:19:@34963.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 73:20:@34957.4]
  assign regs_120_clock = clock; // @[:@34966.4]
  assign regs_120_reset = io_reset; // @[:@34967.4 RegFile.scala 75:16:@34974.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 74:16:@34973.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 77:19:@34977.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 73:20:@34971.4]
  assign regs_121_clock = clock; // @[:@34980.4]
  assign regs_121_reset = io_reset; // @[:@34981.4 RegFile.scala 75:16:@34988.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 74:16:@34987.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 77:19:@34991.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 73:20:@34985.4]
  assign regs_122_clock = clock; // @[:@34994.4]
  assign regs_122_reset = io_reset; // @[:@34995.4 RegFile.scala 75:16:@35002.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 74:16:@35001.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 77:19:@35005.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 73:20:@34999.4]
  assign regs_123_clock = clock; // @[:@35008.4]
  assign regs_123_reset = io_reset; // @[:@35009.4 RegFile.scala 75:16:@35016.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 74:16:@35015.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 77:19:@35019.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 73:20:@35013.4]
  assign regs_124_clock = clock; // @[:@35022.4]
  assign regs_124_reset = io_reset; // @[:@35023.4 RegFile.scala 75:16:@35030.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 74:16:@35029.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 77:19:@35033.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 73:20:@35027.4]
  assign regs_125_clock = clock; // @[:@35036.4]
  assign regs_125_reset = io_reset; // @[:@35037.4 RegFile.scala 75:16:@35044.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 74:16:@35043.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 77:19:@35047.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 73:20:@35041.4]
  assign regs_126_clock = clock; // @[:@35050.4]
  assign regs_126_reset = io_reset; // @[:@35051.4 RegFile.scala 75:16:@35058.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 74:16:@35057.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 77:19:@35061.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 73:20:@35055.4]
  assign regs_127_clock = clock; // @[:@35064.4]
  assign regs_127_reset = io_reset; // @[:@35065.4 RegFile.scala 75:16:@35072.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 74:16:@35071.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 77:19:@35075.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 73:20:@35069.4]
  assign regs_128_clock = clock; // @[:@35078.4]
  assign regs_128_reset = io_reset; // @[:@35079.4 RegFile.scala 75:16:@35086.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 74:16:@35085.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 77:19:@35089.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 73:20:@35083.4]
  assign regs_129_clock = clock; // @[:@35092.4]
  assign regs_129_reset = io_reset; // @[:@35093.4 RegFile.scala 75:16:@35100.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 74:16:@35099.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 77:19:@35103.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 73:20:@35097.4]
  assign regs_130_clock = clock; // @[:@35106.4]
  assign regs_130_reset = io_reset; // @[:@35107.4 RegFile.scala 75:16:@35114.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 74:16:@35113.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 77:19:@35117.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 73:20:@35111.4]
  assign regs_131_clock = clock; // @[:@35120.4]
  assign regs_131_reset = io_reset; // @[:@35121.4 RegFile.scala 75:16:@35128.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 74:16:@35127.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 77:19:@35131.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 73:20:@35125.4]
  assign regs_132_clock = clock; // @[:@35134.4]
  assign regs_132_reset = io_reset; // @[:@35135.4 RegFile.scala 75:16:@35142.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 74:16:@35141.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 77:19:@35145.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 73:20:@35139.4]
  assign regs_133_clock = clock; // @[:@35148.4]
  assign regs_133_reset = io_reset; // @[:@35149.4 RegFile.scala 75:16:@35156.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 74:16:@35155.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 77:19:@35159.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 73:20:@35153.4]
  assign regs_134_clock = clock; // @[:@35162.4]
  assign regs_134_reset = io_reset; // @[:@35163.4 RegFile.scala 75:16:@35170.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 74:16:@35169.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 77:19:@35173.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 73:20:@35167.4]
  assign regs_135_clock = clock; // @[:@35176.4]
  assign regs_135_reset = io_reset; // @[:@35177.4 RegFile.scala 75:16:@35184.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 74:16:@35183.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 77:19:@35187.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 73:20:@35181.4]
  assign regs_136_clock = clock; // @[:@35190.4]
  assign regs_136_reset = io_reset; // @[:@35191.4 RegFile.scala 75:16:@35198.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 74:16:@35197.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 77:19:@35201.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 73:20:@35195.4]
  assign regs_137_clock = clock; // @[:@35204.4]
  assign regs_137_reset = io_reset; // @[:@35205.4 RegFile.scala 75:16:@35212.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 74:16:@35211.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 77:19:@35215.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 73:20:@35209.4]
  assign regs_138_clock = clock; // @[:@35218.4]
  assign regs_138_reset = io_reset; // @[:@35219.4 RegFile.scala 75:16:@35226.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 74:16:@35225.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 77:19:@35229.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 73:20:@35223.4]
  assign regs_139_clock = clock; // @[:@35232.4]
  assign regs_139_reset = io_reset; // @[:@35233.4 RegFile.scala 75:16:@35240.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 74:16:@35239.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 77:19:@35243.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 73:20:@35237.4]
  assign regs_140_clock = clock; // @[:@35246.4]
  assign regs_140_reset = io_reset; // @[:@35247.4 RegFile.scala 75:16:@35254.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 74:16:@35253.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 77:19:@35257.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 73:20:@35251.4]
  assign regs_141_clock = clock; // @[:@35260.4]
  assign regs_141_reset = io_reset; // @[:@35261.4 RegFile.scala 75:16:@35268.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 74:16:@35267.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 77:19:@35271.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 73:20:@35265.4]
  assign regs_142_clock = clock; // @[:@35274.4]
  assign regs_142_reset = io_reset; // @[:@35275.4 RegFile.scala 75:16:@35282.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 74:16:@35281.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 77:19:@35285.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 73:20:@35279.4]
  assign regs_143_clock = clock; // @[:@35288.4]
  assign regs_143_reset = io_reset; // @[:@35289.4 RegFile.scala 75:16:@35296.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 74:16:@35295.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 77:19:@35299.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 73:20:@35293.4]
  assign regs_144_clock = clock; // @[:@35302.4]
  assign regs_144_reset = io_reset; // @[:@35303.4 RegFile.scala 75:16:@35310.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 74:16:@35309.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 77:19:@35313.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 73:20:@35307.4]
  assign regs_145_clock = clock; // @[:@35316.4]
  assign regs_145_reset = io_reset; // @[:@35317.4 RegFile.scala 75:16:@35324.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 74:16:@35323.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 77:19:@35327.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 73:20:@35321.4]
  assign regs_146_clock = clock; // @[:@35330.4]
  assign regs_146_reset = io_reset; // @[:@35331.4 RegFile.scala 75:16:@35338.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 74:16:@35337.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 77:19:@35341.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 73:20:@35335.4]
  assign regs_147_clock = clock; // @[:@35344.4]
  assign regs_147_reset = io_reset; // @[:@35345.4 RegFile.scala 75:16:@35352.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 74:16:@35351.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 77:19:@35355.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 73:20:@35349.4]
  assign regs_148_clock = clock; // @[:@35358.4]
  assign regs_148_reset = io_reset; // @[:@35359.4 RegFile.scala 75:16:@35366.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 74:16:@35365.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 77:19:@35369.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 73:20:@35363.4]
  assign regs_149_clock = clock; // @[:@35372.4]
  assign regs_149_reset = io_reset; // @[:@35373.4 RegFile.scala 75:16:@35380.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 74:16:@35379.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 77:19:@35383.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 73:20:@35377.4]
  assign regs_150_clock = clock; // @[:@35386.4]
  assign regs_150_reset = io_reset; // @[:@35387.4 RegFile.scala 75:16:@35394.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 74:16:@35393.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 77:19:@35397.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 73:20:@35391.4]
  assign regs_151_clock = clock; // @[:@35400.4]
  assign regs_151_reset = io_reset; // @[:@35401.4 RegFile.scala 75:16:@35408.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 74:16:@35407.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 77:19:@35411.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 73:20:@35405.4]
  assign regs_152_clock = clock; // @[:@35414.4]
  assign regs_152_reset = io_reset; // @[:@35415.4 RegFile.scala 75:16:@35422.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 74:16:@35421.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 77:19:@35425.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 73:20:@35419.4]
  assign regs_153_clock = clock; // @[:@35428.4]
  assign regs_153_reset = io_reset; // @[:@35429.4 RegFile.scala 75:16:@35436.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 74:16:@35435.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 77:19:@35439.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 73:20:@35433.4]
  assign regs_154_clock = clock; // @[:@35442.4]
  assign regs_154_reset = io_reset; // @[:@35443.4 RegFile.scala 75:16:@35450.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 74:16:@35449.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 77:19:@35453.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 73:20:@35447.4]
  assign regs_155_clock = clock; // @[:@35456.4]
  assign regs_155_reset = io_reset; // @[:@35457.4 RegFile.scala 75:16:@35464.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 74:16:@35463.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 77:19:@35467.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 73:20:@35461.4]
  assign regs_156_clock = clock; // @[:@35470.4]
  assign regs_156_reset = io_reset; // @[:@35471.4 RegFile.scala 75:16:@35478.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 74:16:@35477.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 77:19:@35481.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 73:20:@35475.4]
  assign regs_157_clock = clock; // @[:@35484.4]
  assign regs_157_reset = io_reset; // @[:@35485.4 RegFile.scala 75:16:@35492.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 74:16:@35491.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 77:19:@35495.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 73:20:@35489.4]
  assign regs_158_clock = clock; // @[:@35498.4]
  assign regs_158_reset = io_reset; // @[:@35499.4 RegFile.scala 75:16:@35506.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 74:16:@35505.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 77:19:@35509.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 73:20:@35503.4]
  assign regs_159_clock = clock; // @[:@35512.4]
  assign regs_159_reset = io_reset; // @[:@35513.4 RegFile.scala 75:16:@35520.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 74:16:@35519.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 77:19:@35523.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 73:20:@35517.4]
  assign regs_160_clock = clock; // @[:@35526.4]
  assign regs_160_reset = io_reset; // @[:@35527.4 RegFile.scala 75:16:@35534.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 74:16:@35533.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 77:19:@35537.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 73:20:@35531.4]
  assign regs_161_clock = clock; // @[:@35540.4]
  assign regs_161_reset = io_reset; // @[:@35541.4 RegFile.scala 75:16:@35548.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 74:16:@35547.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 77:19:@35551.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 73:20:@35545.4]
  assign regs_162_clock = clock; // @[:@35554.4]
  assign regs_162_reset = io_reset; // @[:@35555.4 RegFile.scala 75:16:@35562.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 74:16:@35561.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 77:19:@35565.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 73:20:@35559.4]
  assign regs_163_clock = clock; // @[:@35568.4]
  assign regs_163_reset = io_reset; // @[:@35569.4 RegFile.scala 75:16:@35576.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 74:16:@35575.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 77:19:@35579.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 73:20:@35573.4]
  assign regs_164_clock = clock; // @[:@35582.4]
  assign regs_164_reset = io_reset; // @[:@35583.4 RegFile.scala 75:16:@35590.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 74:16:@35589.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 77:19:@35593.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 73:20:@35587.4]
  assign regs_165_clock = clock; // @[:@35596.4]
  assign regs_165_reset = io_reset; // @[:@35597.4 RegFile.scala 75:16:@35604.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 74:16:@35603.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 77:19:@35607.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 73:20:@35601.4]
  assign regs_166_clock = clock; // @[:@35610.4]
  assign regs_166_reset = io_reset; // @[:@35611.4 RegFile.scala 75:16:@35618.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 74:16:@35617.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 77:19:@35621.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 73:20:@35615.4]
  assign regs_167_clock = clock; // @[:@35624.4]
  assign regs_167_reset = io_reset; // @[:@35625.4 RegFile.scala 75:16:@35632.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 74:16:@35631.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 77:19:@35635.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 73:20:@35629.4]
  assign regs_168_clock = clock; // @[:@35638.4]
  assign regs_168_reset = io_reset; // @[:@35639.4 RegFile.scala 75:16:@35646.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 74:16:@35645.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 77:19:@35649.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 73:20:@35643.4]
  assign regs_169_clock = clock; // @[:@35652.4]
  assign regs_169_reset = io_reset; // @[:@35653.4 RegFile.scala 75:16:@35660.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 74:16:@35659.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 77:19:@35663.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 73:20:@35657.4]
  assign regs_170_clock = clock; // @[:@35666.4]
  assign regs_170_reset = io_reset; // @[:@35667.4 RegFile.scala 75:16:@35674.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 74:16:@35673.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 77:19:@35677.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 73:20:@35671.4]
  assign regs_171_clock = clock; // @[:@35680.4]
  assign regs_171_reset = io_reset; // @[:@35681.4 RegFile.scala 75:16:@35688.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 74:16:@35687.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 77:19:@35691.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 73:20:@35685.4]
  assign regs_172_clock = clock; // @[:@35694.4]
  assign regs_172_reset = io_reset; // @[:@35695.4 RegFile.scala 75:16:@35702.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 74:16:@35701.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 77:19:@35705.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 73:20:@35699.4]
  assign regs_173_clock = clock; // @[:@35708.4]
  assign regs_173_reset = io_reset; // @[:@35709.4 RegFile.scala 75:16:@35716.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 74:16:@35715.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 77:19:@35719.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 73:20:@35713.4]
  assign regs_174_clock = clock; // @[:@35722.4]
  assign regs_174_reset = io_reset; // @[:@35723.4 RegFile.scala 75:16:@35730.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 74:16:@35729.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 77:19:@35733.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 73:20:@35727.4]
  assign regs_175_clock = clock; // @[:@35736.4]
  assign regs_175_reset = io_reset; // @[:@35737.4 RegFile.scala 75:16:@35744.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 74:16:@35743.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 77:19:@35747.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 73:20:@35741.4]
  assign regs_176_clock = clock; // @[:@35750.4]
  assign regs_176_reset = io_reset; // @[:@35751.4 RegFile.scala 75:16:@35758.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 74:16:@35757.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 77:19:@35761.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 73:20:@35755.4]
  assign regs_177_clock = clock; // @[:@35764.4]
  assign regs_177_reset = io_reset; // @[:@35765.4 RegFile.scala 75:16:@35772.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 74:16:@35771.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 77:19:@35775.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 73:20:@35769.4]
  assign regs_178_clock = clock; // @[:@35778.4]
  assign regs_178_reset = io_reset; // @[:@35779.4 RegFile.scala 75:16:@35786.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 74:16:@35785.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 77:19:@35789.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 73:20:@35783.4]
  assign regs_179_clock = clock; // @[:@35792.4]
  assign regs_179_reset = io_reset; // @[:@35793.4 RegFile.scala 75:16:@35800.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 74:16:@35799.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 77:19:@35803.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 73:20:@35797.4]
  assign regs_180_clock = clock; // @[:@35806.4]
  assign regs_180_reset = io_reset; // @[:@35807.4 RegFile.scala 75:16:@35814.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 74:16:@35813.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 77:19:@35817.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 73:20:@35811.4]
  assign regs_181_clock = clock; // @[:@35820.4]
  assign regs_181_reset = io_reset; // @[:@35821.4 RegFile.scala 75:16:@35828.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 74:16:@35827.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 77:19:@35831.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 73:20:@35825.4]
  assign regs_182_clock = clock; // @[:@35834.4]
  assign regs_182_reset = io_reset; // @[:@35835.4 RegFile.scala 75:16:@35842.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 74:16:@35841.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 77:19:@35845.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 73:20:@35839.4]
  assign regs_183_clock = clock; // @[:@35848.4]
  assign regs_183_reset = io_reset; // @[:@35849.4 RegFile.scala 75:16:@35856.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 74:16:@35855.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 77:19:@35859.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 73:20:@35853.4]
  assign regs_184_clock = clock; // @[:@35862.4]
  assign regs_184_reset = io_reset; // @[:@35863.4 RegFile.scala 75:16:@35870.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 74:16:@35869.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 77:19:@35873.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 73:20:@35867.4]
  assign regs_185_clock = clock; // @[:@35876.4]
  assign regs_185_reset = io_reset; // @[:@35877.4 RegFile.scala 75:16:@35884.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 74:16:@35883.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 77:19:@35887.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 73:20:@35881.4]
  assign regs_186_clock = clock; // @[:@35890.4]
  assign regs_186_reset = io_reset; // @[:@35891.4 RegFile.scala 75:16:@35898.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 74:16:@35897.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 77:19:@35901.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 73:20:@35895.4]
  assign regs_187_clock = clock; // @[:@35904.4]
  assign regs_187_reset = io_reset; // @[:@35905.4 RegFile.scala 75:16:@35912.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 74:16:@35911.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 77:19:@35915.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 73:20:@35909.4]
  assign regs_188_clock = clock; // @[:@35918.4]
  assign regs_188_reset = io_reset; // @[:@35919.4 RegFile.scala 75:16:@35926.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 74:16:@35925.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 77:19:@35929.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 73:20:@35923.4]
  assign regs_189_clock = clock; // @[:@35932.4]
  assign regs_189_reset = io_reset; // @[:@35933.4 RegFile.scala 75:16:@35940.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 74:16:@35939.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 77:19:@35943.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 73:20:@35937.4]
  assign regs_190_clock = clock; // @[:@35946.4]
  assign regs_190_reset = io_reset; // @[:@35947.4 RegFile.scala 75:16:@35954.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 74:16:@35953.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 77:19:@35957.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 73:20:@35951.4]
  assign regs_191_clock = clock; // @[:@35960.4]
  assign regs_191_reset = io_reset; // @[:@35961.4 RegFile.scala 75:16:@35968.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 74:16:@35967.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 77:19:@35971.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 73:20:@35965.4]
  assign regs_192_clock = clock; // @[:@35974.4]
  assign regs_192_reset = io_reset; // @[:@35975.4 RegFile.scala 75:16:@35982.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 74:16:@35981.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 77:19:@35985.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 73:20:@35979.4]
  assign regs_193_clock = clock; // @[:@35988.4]
  assign regs_193_reset = io_reset; // @[:@35989.4 RegFile.scala 75:16:@35996.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 74:16:@35995.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 77:19:@35999.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 73:20:@35993.4]
  assign regs_194_clock = clock; // @[:@36002.4]
  assign regs_194_reset = io_reset; // @[:@36003.4 RegFile.scala 75:16:@36010.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 74:16:@36009.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 77:19:@36013.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 73:20:@36007.4]
  assign regs_195_clock = clock; // @[:@36016.4]
  assign regs_195_reset = io_reset; // @[:@36017.4 RegFile.scala 75:16:@36024.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 74:16:@36023.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 77:19:@36027.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 73:20:@36021.4]
  assign regs_196_clock = clock; // @[:@36030.4]
  assign regs_196_reset = io_reset; // @[:@36031.4 RegFile.scala 75:16:@36038.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 74:16:@36037.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 77:19:@36041.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 73:20:@36035.4]
  assign regs_197_clock = clock; // @[:@36044.4]
  assign regs_197_reset = io_reset; // @[:@36045.4 RegFile.scala 75:16:@36052.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 74:16:@36051.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 77:19:@36055.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 73:20:@36049.4]
  assign regs_198_clock = clock; // @[:@36058.4]
  assign regs_198_reset = io_reset; // @[:@36059.4 RegFile.scala 75:16:@36066.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 74:16:@36065.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 77:19:@36069.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 73:20:@36063.4]
  assign regs_199_clock = clock; // @[:@36072.4]
  assign regs_199_reset = io_reset; // @[:@36073.4 RegFile.scala 75:16:@36080.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 74:16:@36079.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 77:19:@36083.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 73:20:@36077.4]
  assign regs_200_clock = clock; // @[:@36086.4]
  assign regs_200_reset = io_reset; // @[:@36087.4 RegFile.scala 75:16:@36094.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 74:16:@36093.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 77:19:@36097.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 73:20:@36091.4]
  assign regs_201_clock = clock; // @[:@36100.4]
  assign regs_201_reset = io_reset; // @[:@36101.4 RegFile.scala 75:16:@36108.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 74:16:@36107.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 77:19:@36111.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 73:20:@36105.4]
  assign regs_202_clock = clock; // @[:@36114.4]
  assign regs_202_reset = io_reset; // @[:@36115.4 RegFile.scala 75:16:@36122.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 74:16:@36121.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 77:19:@36125.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 73:20:@36119.4]
  assign regs_203_clock = clock; // @[:@36128.4]
  assign regs_203_reset = io_reset; // @[:@36129.4 RegFile.scala 75:16:@36136.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 74:16:@36135.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 77:19:@36139.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 73:20:@36133.4]
  assign regs_204_clock = clock; // @[:@36142.4]
  assign regs_204_reset = io_reset; // @[:@36143.4 RegFile.scala 75:16:@36150.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 74:16:@36149.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 77:19:@36153.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 73:20:@36147.4]
  assign regs_205_clock = clock; // @[:@36156.4]
  assign regs_205_reset = io_reset; // @[:@36157.4 RegFile.scala 75:16:@36164.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 74:16:@36163.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 77:19:@36167.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 73:20:@36161.4]
  assign regs_206_clock = clock; // @[:@36170.4]
  assign regs_206_reset = io_reset; // @[:@36171.4 RegFile.scala 75:16:@36178.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 74:16:@36177.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 77:19:@36181.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 73:20:@36175.4]
  assign regs_207_clock = clock; // @[:@36184.4]
  assign regs_207_reset = io_reset; // @[:@36185.4 RegFile.scala 75:16:@36192.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 74:16:@36191.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 77:19:@36195.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 73:20:@36189.4]
  assign regs_208_clock = clock; // @[:@36198.4]
  assign regs_208_reset = io_reset; // @[:@36199.4 RegFile.scala 75:16:@36206.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 74:16:@36205.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 77:19:@36209.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 73:20:@36203.4]
  assign regs_209_clock = clock; // @[:@36212.4]
  assign regs_209_reset = io_reset; // @[:@36213.4 RegFile.scala 75:16:@36220.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 74:16:@36219.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 77:19:@36223.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 73:20:@36217.4]
  assign regs_210_clock = clock; // @[:@36226.4]
  assign regs_210_reset = io_reset; // @[:@36227.4 RegFile.scala 75:16:@36234.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 74:16:@36233.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 77:19:@36237.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 73:20:@36231.4]
  assign regs_211_clock = clock; // @[:@36240.4]
  assign regs_211_reset = io_reset; // @[:@36241.4 RegFile.scala 75:16:@36248.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 74:16:@36247.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 77:19:@36251.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 73:20:@36245.4]
  assign regs_212_clock = clock; // @[:@36254.4]
  assign regs_212_reset = io_reset; // @[:@36255.4 RegFile.scala 75:16:@36262.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 74:16:@36261.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 77:19:@36265.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 73:20:@36259.4]
  assign regs_213_clock = clock; // @[:@36268.4]
  assign regs_213_reset = io_reset; // @[:@36269.4 RegFile.scala 75:16:@36276.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 74:16:@36275.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 77:19:@36279.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 73:20:@36273.4]
  assign regs_214_clock = clock; // @[:@36282.4]
  assign regs_214_reset = io_reset; // @[:@36283.4 RegFile.scala 75:16:@36290.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 74:16:@36289.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 77:19:@36293.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 73:20:@36287.4]
  assign regs_215_clock = clock; // @[:@36296.4]
  assign regs_215_reset = io_reset; // @[:@36297.4 RegFile.scala 75:16:@36304.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 74:16:@36303.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 77:19:@36307.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 73:20:@36301.4]
  assign regs_216_clock = clock; // @[:@36310.4]
  assign regs_216_reset = io_reset; // @[:@36311.4 RegFile.scala 75:16:@36318.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 74:16:@36317.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 77:19:@36321.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 73:20:@36315.4]
  assign regs_217_clock = clock; // @[:@36324.4]
  assign regs_217_reset = io_reset; // @[:@36325.4 RegFile.scala 75:16:@36332.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 74:16:@36331.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 77:19:@36335.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 73:20:@36329.4]
  assign regs_218_clock = clock; // @[:@36338.4]
  assign regs_218_reset = io_reset; // @[:@36339.4 RegFile.scala 75:16:@36346.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 74:16:@36345.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 77:19:@36349.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 73:20:@36343.4]
  assign regs_219_clock = clock; // @[:@36352.4]
  assign regs_219_reset = io_reset; // @[:@36353.4 RegFile.scala 75:16:@36360.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 74:16:@36359.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 77:19:@36363.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 73:20:@36357.4]
  assign regs_220_clock = clock; // @[:@36366.4]
  assign regs_220_reset = io_reset; // @[:@36367.4 RegFile.scala 75:16:@36374.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 74:16:@36373.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 77:19:@36377.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 73:20:@36371.4]
  assign regs_221_clock = clock; // @[:@36380.4]
  assign regs_221_reset = io_reset; // @[:@36381.4 RegFile.scala 75:16:@36388.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 74:16:@36387.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 77:19:@36391.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 73:20:@36385.4]
  assign regs_222_clock = clock; // @[:@36394.4]
  assign regs_222_reset = io_reset; // @[:@36395.4 RegFile.scala 75:16:@36402.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 74:16:@36401.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 77:19:@36405.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 73:20:@36399.4]
  assign regs_223_clock = clock; // @[:@36408.4]
  assign regs_223_reset = io_reset; // @[:@36409.4 RegFile.scala 75:16:@36416.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 74:16:@36415.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 77:19:@36419.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 73:20:@36413.4]
  assign regs_224_clock = clock; // @[:@36422.4]
  assign regs_224_reset = io_reset; // @[:@36423.4 RegFile.scala 75:16:@36430.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 74:16:@36429.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 77:19:@36433.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 73:20:@36427.4]
  assign regs_225_clock = clock; // @[:@36436.4]
  assign regs_225_reset = io_reset; // @[:@36437.4 RegFile.scala 75:16:@36444.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 74:16:@36443.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 77:19:@36447.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 73:20:@36441.4]
  assign regs_226_clock = clock; // @[:@36450.4]
  assign regs_226_reset = io_reset; // @[:@36451.4 RegFile.scala 75:16:@36458.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 74:16:@36457.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 77:19:@36461.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 73:20:@36455.4]
  assign regs_227_clock = clock; // @[:@36464.4]
  assign regs_227_reset = io_reset; // @[:@36465.4 RegFile.scala 75:16:@36472.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 74:16:@36471.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 77:19:@36475.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 73:20:@36469.4]
  assign regs_228_clock = clock; // @[:@36478.4]
  assign regs_228_reset = io_reset; // @[:@36479.4 RegFile.scala 75:16:@36486.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 74:16:@36485.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 77:19:@36489.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 73:20:@36483.4]
  assign regs_229_clock = clock; // @[:@36492.4]
  assign regs_229_reset = io_reset; // @[:@36493.4 RegFile.scala 75:16:@36500.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 74:16:@36499.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 77:19:@36503.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 73:20:@36497.4]
  assign regs_230_clock = clock; // @[:@36506.4]
  assign regs_230_reset = io_reset; // @[:@36507.4 RegFile.scala 75:16:@36514.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 74:16:@36513.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 77:19:@36517.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 73:20:@36511.4]
  assign regs_231_clock = clock; // @[:@36520.4]
  assign regs_231_reset = io_reset; // @[:@36521.4 RegFile.scala 75:16:@36528.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 74:16:@36527.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 77:19:@36531.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 73:20:@36525.4]
  assign regs_232_clock = clock; // @[:@36534.4]
  assign regs_232_reset = io_reset; // @[:@36535.4 RegFile.scala 75:16:@36542.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 74:16:@36541.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 77:19:@36545.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 73:20:@36539.4]
  assign regs_233_clock = clock; // @[:@36548.4]
  assign regs_233_reset = io_reset; // @[:@36549.4 RegFile.scala 75:16:@36556.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 74:16:@36555.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 77:19:@36559.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 73:20:@36553.4]
  assign regs_234_clock = clock; // @[:@36562.4]
  assign regs_234_reset = io_reset; // @[:@36563.4 RegFile.scala 75:16:@36570.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 74:16:@36569.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 77:19:@36573.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 73:20:@36567.4]
  assign regs_235_clock = clock; // @[:@36576.4]
  assign regs_235_reset = io_reset; // @[:@36577.4 RegFile.scala 75:16:@36584.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 74:16:@36583.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 77:19:@36587.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 73:20:@36581.4]
  assign regs_236_clock = clock; // @[:@36590.4]
  assign regs_236_reset = io_reset; // @[:@36591.4 RegFile.scala 75:16:@36598.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 74:16:@36597.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 77:19:@36601.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 73:20:@36595.4]
  assign regs_237_clock = clock; // @[:@36604.4]
  assign regs_237_reset = io_reset; // @[:@36605.4 RegFile.scala 75:16:@36612.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 74:16:@36611.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 77:19:@36615.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 73:20:@36609.4]
  assign regs_238_clock = clock; // @[:@36618.4]
  assign regs_238_reset = io_reset; // @[:@36619.4 RegFile.scala 75:16:@36626.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 74:16:@36625.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 77:19:@36629.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 73:20:@36623.4]
  assign regs_239_clock = clock; // @[:@36632.4]
  assign regs_239_reset = io_reset; // @[:@36633.4 RegFile.scala 75:16:@36640.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 74:16:@36639.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 77:19:@36643.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 73:20:@36637.4]
  assign regs_240_clock = clock; // @[:@36646.4]
  assign regs_240_reset = io_reset; // @[:@36647.4 RegFile.scala 75:16:@36654.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 74:16:@36653.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 77:19:@36657.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 73:20:@36651.4]
  assign regs_241_clock = clock; // @[:@36660.4]
  assign regs_241_reset = io_reset; // @[:@36661.4 RegFile.scala 75:16:@36668.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 74:16:@36667.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 77:19:@36671.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 73:20:@36665.4]
  assign regs_242_clock = clock; // @[:@36674.4]
  assign regs_242_reset = io_reset; // @[:@36675.4 RegFile.scala 75:16:@36682.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 74:16:@36681.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 77:19:@36685.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 73:20:@36679.4]
  assign regs_243_clock = clock; // @[:@36688.4]
  assign regs_243_reset = io_reset; // @[:@36689.4 RegFile.scala 75:16:@36696.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 74:16:@36695.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 77:19:@36699.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 73:20:@36693.4]
  assign regs_244_clock = clock; // @[:@36702.4]
  assign regs_244_reset = io_reset; // @[:@36703.4 RegFile.scala 75:16:@36710.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 74:16:@36709.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 77:19:@36713.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 73:20:@36707.4]
  assign regs_245_clock = clock; // @[:@36716.4]
  assign regs_245_reset = io_reset; // @[:@36717.4 RegFile.scala 75:16:@36724.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 74:16:@36723.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 77:19:@36727.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 73:20:@36721.4]
  assign regs_246_clock = clock; // @[:@36730.4]
  assign regs_246_reset = io_reset; // @[:@36731.4 RegFile.scala 75:16:@36738.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 74:16:@36737.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 77:19:@36741.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 73:20:@36735.4]
  assign regs_247_clock = clock; // @[:@36744.4]
  assign regs_247_reset = io_reset; // @[:@36745.4 RegFile.scala 75:16:@36752.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 74:16:@36751.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 77:19:@36755.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 73:20:@36749.4]
  assign regs_248_clock = clock; // @[:@36758.4]
  assign regs_248_reset = io_reset; // @[:@36759.4 RegFile.scala 75:16:@36766.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 74:16:@36765.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 77:19:@36769.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 73:20:@36763.4]
  assign regs_249_clock = clock; // @[:@36772.4]
  assign regs_249_reset = io_reset; // @[:@36773.4 RegFile.scala 75:16:@36780.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 74:16:@36779.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 77:19:@36783.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 73:20:@36777.4]
  assign regs_250_clock = clock; // @[:@36786.4]
  assign regs_250_reset = io_reset; // @[:@36787.4 RegFile.scala 75:16:@36794.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 74:16:@36793.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 77:19:@36797.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 73:20:@36791.4]
  assign regs_251_clock = clock; // @[:@36800.4]
  assign regs_251_reset = io_reset; // @[:@36801.4 RegFile.scala 75:16:@36808.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 74:16:@36807.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 77:19:@36811.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 73:20:@36805.4]
  assign regs_252_clock = clock; // @[:@36814.4]
  assign regs_252_reset = io_reset; // @[:@36815.4 RegFile.scala 75:16:@36822.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 74:16:@36821.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 77:19:@36825.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 73:20:@36819.4]
  assign regs_253_clock = clock; // @[:@36828.4]
  assign regs_253_reset = io_reset; // @[:@36829.4 RegFile.scala 75:16:@36836.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 74:16:@36835.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 77:19:@36839.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 73:20:@36833.4]
  assign regs_254_clock = clock; // @[:@36842.4]
  assign regs_254_reset = io_reset; // @[:@36843.4 RegFile.scala 75:16:@36850.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 74:16:@36849.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 77:19:@36853.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 73:20:@36847.4]
  assign regs_255_clock = clock; // @[:@36856.4]
  assign regs_255_reset = io_reset; // @[:@36857.4 RegFile.scala 75:16:@36864.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 74:16:@36863.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 77:19:@36867.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 73:20:@36861.4]
  assign regs_256_clock = clock; // @[:@36870.4]
  assign regs_256_reset = io_reset; // @[:@36871.4 RegFile.scala 75:16:@36878.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 74:16:@36877.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 77:19:@36881.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 73:20:@36875.4]
  assign regs_257_clock = clock; // @[:@36884.4]
  assign regs_257_reset = io_reset; // @[:@36885.4 RegFile.scala 75:16:@36892.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 74:16:@36891.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 77:19:@36895.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 73:20:@36889.4]
  assign regs_258_clock = clock; // @[:@36898.4]
  assign regs_258_reset = io_reset; // @[:@36899.4 RegFile.scala 75:16:@36906.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 74:16:@36905.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 77:19:@36909.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 73:20:@36903.4]
  assign regs_259_clock = clock; // @[:@36912.4]
  assign regs_259_reset = io_reset; // @[:@36913.4 RegFile.scala 75:16:@36920.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 74:16:@36919.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 77:19:@36923.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 73:20:@36917.4]
  assign regs_260_clock = clock; // @[:@36926.4]
  assign regs_260_reset = io_reset; // @[:@36927.4 RegFile.scala 75:16:@36934.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 74:16:@36933.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 77:19:@36937.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 73:20:@36931.4]
  assign regs_261_clock = clock; // @[:@36940.4]
  assign regs_261_reset = io_reset; // @[:@36941.4 RegFile.scala 75:16:@36948.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 74:16:@36947.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 77:19:@36951.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 73:20:@36945.4]
  assign regs_262_clock = clock; // @[:@36954.4]
  assign regs_262_reset = io_reset; // @[:@36955.4 RegFile.scala 75:16:@36962.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 74:16:@36961.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 77:19:@36965.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 73:20:@36959.4]
  assign regs_263_clock = clock; // @[:@36968.4]
  assign regs_263_reset = io_reset; // @[:@36969.4 RegFile.scala 75:16:@36976.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 74:16:@36975.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 77:19:@36979.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 73:20:@36973.4]
  assign regs_264_clock = clock; // @[:@36982.4]
  assign regs_264_reset = io_reset; // @[:@36983.4 RegFile.scala 75:16:@36990.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 74:16:@36989.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 77:19:@36993.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 73:20:@36987.4]
  assign regs_265_clock = clock; // @[:@36996.4]
  assign regs_265_reset = io_reset; // @[:@36997.4 RegFile.scala 75:16:@37004.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 74:16:@37003.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 77:19:@37007.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 73:20:@37001.4]
  assign regs_266_clock = clock; // @[:@37010.4]
  assign regs_266_reset = io_reset; // @[:@37011.4 RegFile.scala 75:16:@37018.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 74:16:@37017.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 77:19:@37021.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 73:20:@37015.4]
  assign regs_267_clock = clock; // @[:@37024.4]
  assign regs_267_reset = io_reset; // @[:@37025.4 RegFile.scala 75:16:@37032.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 74:16:@37031.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 77:19:@37035.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 73:20:@37029.4]
  assign regs_268_clock = clock; // @[:@37038.4]
  assign regs_268_reset = io_reset; // @[:@37039.4 RegFile.scala 75:16:@37046.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 74:16:@37045.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 77:19:@37049.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 73:20:@37043.4]
  assign regs_269_clock = clock; // @[:@37052.4]
  assign regs_269_reset = io_reset; // @[:@37053.4 RegFile.scala 75:16:@37060.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 74:16:@37059.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 77:19:@37063.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 73:20:@37057.4]
  assign regs_270_clock = clock; // @[:@37066.4]
  assign regs_270_reset = io_reset; // @[:@37067.4 RegFile.scala 75:16:@37074.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 74:16:@37073.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 77:19:@37077.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 73:20:@37071.4]
  assign regs_271_clock = clock; // @[:@37080.4]
  assign regs_271_reset = io_reset; // @[:@37081.4 RegFile.scala 75:16:@37088.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 74:16:@37087.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 77:19:@37091.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 73:20:@37085.4]
  assign regs_272_clock = clock; // @[:@37094.4]
  assign regs_272_reset = io_reset; // @[:@37095.4 RegFile.scala 75:16:@37102.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 74:16:@37101.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 77:19:@37105.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 73:20:@37099.4]
  assign regs_273_clock = clock; // @[:@37108.4]
  assign regs_273_reset = io_reset; // @[:@37109.4 RegFile.scala 75:16:@37116.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 74:16:@37115.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 77:19:@37119.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 73:20:@37113.4]
  assign regs_274_clock = clock; // @[:@37122.4]
  assign regs_274_reset = io_reset; // @[:@37123.4 RegFile.scala 75:16:@37130.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 74:16:@37129.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 77:19:@37133.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 73:20:@37127.4]
  assign regs_275_clock = clock; // @[:@37136.4]
  assign regs_275_reset = io_reset; // @[:@37137.4 RegFile.scala 75:16:@37144.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 74:16:@37143.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 77:19:@37147.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 73:20:@37141.4]
  assign regs_276_clock = clock; // @[:@37150.4]
  assign regs_276_reset = io_reset; // @[:@37151.4 RegFile.scala 75:16:@37158.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 74:16:@37157.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 77:19:@37161.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 73:20:@37155.4]
  assign regs_277_clock = clock; // @[:@37164.4]
  assign regs_277_reset = io_reset; // @[:@37165.4 RegFile.scala 75:16:@37172.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 74:16:@37171.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 77:19:@37175.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 73:20:@37169.4]
  assign regs_278_clock = clock; // @[:@37178.4]
  assign regs_278_reset = io_reset; // @[:@37179.4 RegFile.scala 75:16:@37186.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 74:16:@37185.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 77:19:@37189.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 73:20:@37183.4]
  assign regs_279_clock = clock; // @[:@37192.4]
  assign regs_279_reset = io_reset; // @[:@37193.4 RegFile.scala 75:16:@37200.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 74:16:@37199.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 77:19:@37203.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 73:20:@37197.4]
  assign regs_280_clock = clock; // @[:@37206.4]
  assign regs_280_reset = io_reset; // @[:@37207.4 RegFile.scala 75:16:@37214.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 74:16:@37213.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 77:19:@37217.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 73:20:@37211.4]
  assign regs_281_clock = clock; // @[:@37220.4]
  assign regs_281_reset = io_reset; // @[:@37221.4 RegFile.scala 75:16:@37228.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 74:16:@37227.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 77:19:@37231.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 73:20:@37225.4]
  assign regs_282_clock = clock; // @[:@37234.4]
  assign regs_282_reset = io_reset; // @[:@37235.4 RegFile.scala 75:16:@37242.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 74:16:@37241.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 77:19:@37245.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 73:20:@37239.4]
  assign regs_283_clock = clock; // @[:@37248.4]
  assign regs_283_reset = io_reset; // @[:@37249.4 RegFile.scala 75:16:@37256.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 74:16:@37255.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 77:19:@37259.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 73:20:@37253.4]
  assign regs_284_clock = clock; // @[:@37262.4]
  assign regs_284_reset = io_reset; // @[:@37263.4 RegFile.scala 75:16:@37270.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 74:16:@37269.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 77:19:@37273.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 73:20:@37267.4]
  assign regs_285_clock = clock; // @[:@37276.4]
  assign regs_285_reset = io_reset; // @[:@37277.4 RegFile.scala 75:16:@37284.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 74:16:@37283.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 77:19:@37287.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 73:20:@37281.4]
  assign regs_286_clock = clock; // @[:@37290.4]
  assign regs_286_reset = io_reset; // @[:@37291.4 RegFile.scala 75:16:@37298.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 74:16:@37297.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 77:19:@37301.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 73:20:@37295.4]
  assign regs_287_clock = clock; // @[:@37304.4]
  assign regs_287_reset = io_reset; // @[:@37305.4 RegFile.scala 75:16:@37312.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 74:16:@37311.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 77:19:@37315.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 73:20:@37309.4]
  assign regs_288_clock = clock; // @[:@37318.4]
  assign regs_288_reset = io_reset; // @[:@37319.4 RegFile.scala 75:16:@37326.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 74:16:@37325.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 77:19:@37329.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 73:20:@37323.4]
  assign regs_289_clock = clock; // @[:@37332.4]
  assign regs_289_reset = io_reset; // @[:@37333.4 RegFile.scala 75:16:@37340.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 74:16:@37339.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 77:19:@37343.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 73:20:@37337.4]
  assign regs_290_clock = clock; // @[:@37346.4]
  assign regs_290_reset = io_reset; // @[:@37347.4 RegFile.scala 75:16:@37354.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 74:16:@37353.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 77:19:@37357.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 73:20:@37351.4]
  assign regs_291_clock = clock; // @[:@37360.4]
  assign regs_291_reset = io_reset; // @[:@37361.4 RegFile.scala 75:16:@37368.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 74:16:@37367.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 77:19:@37371.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 73:20:@37365.4]
  assign regs_292_clock = clock; // @[:@37374.4]
  assign regs_292_reset = io_reset; // @[:@37375.4 RegFile.scala 75:16:@37382.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 74:16:@37381.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 77:19:@37385.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 73:20:@37379.4]
  assign regs_293_clock = clock; // @[:@37388.4]
  assign regs_293_reset = io_reset; // @[:@37389.4 RegFile.scala 75:16:@37396.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 74:16:@37395.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 77:19:@37399.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 73:20:@37393.4]
  assign regs_294_clock = clock; // @[:@37402.4]
  assign regs_294_reset = io_reset; // @[:@37403.4 RegFile.scala 75:16:@37410.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 74:16:@37409.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 77:19:@37413.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 73:20:@37407.4]
  assign regs_295_clock = clock; // @[:@37416.4]
  assign regs_295_reset = io_reset; // @[:@37417.4 RegFile.scala 75:16:@37424.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 74:16:@37423.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 77:19:@37427.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 73:20:@37421.4]
  assign regs_296_clock = clock; // @[:@37430.4]
  assign regs_296_reset = io_reset; // @[:@37431.4 RegFile.scala 75:16:@37438.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 74:16:@37437.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 77:19:@37441.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 73:20:@37435.4]
  assign regs_297_clock = clock; // @[:@37444.4]
  assign regs_297_reset = io_reset; // @[:@37445.4 RegFile.scala 75:16:@37452.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 74:16:@37451.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 77:19:@37455.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 73:20:@37449.4]
  assign regs_298_clock = clock; // @[:@37458.4]
  assign regs_298_reset = io_reset; // @[:@37459.4 RegFile.scala 75:16:@37466.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 74:16:@37465.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 77:19:@37469.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 73:20:@37463.4]
  assign regs_299_clock = clock; // @[:@37472.4]
  assign regs_299_reset = io_reset; // @[:@37473.4 RegFile.scala 75:16:@37480.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 74:16:@37479.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 77:19:@37483.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 73:20:@37477.4]
  assign regs_300_clock = clock; // @[:@37486.4]
  assign regs_300_reset = io_reset; // @[:@37487.4 RegFile.scala 75:16:@37494.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 74:16:@37493.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 77:19:@37497.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 73:20:@37491.4]
  assign regs_301_clock = clock; // @[:@37500.4]
  assign regs_301_reset = io_reset; // @[:@37501.4 RegFile.scala 75:16:@37508.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 74:16:@37507.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 77:19:@37511.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 73:20:@37505.4]
  assign regs_302_clock = clock; // @[:@37514.4]
  assign regs_302_reset = io_reset; // @[:@37515.4 RegFile.scala 75:16:@37522.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 74:16:@37521.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 77:19:@37525.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 73:20:@37519.4]
  assign regs_303_clock = clock; // @[:@37528.4]
  assign regs_303_reset = io_reset; // @[:@37529.4 RegFile.scala 75:16:@37536.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 74:16:@37535.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 77:19:@37539.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 73:20:@37533.4]
  assign regs_304_clock = clock; // @[:@37542.4]
  assign regs_304_reset = io_reset; // @[:@37543.4 RegFile.scala 75:16:@37550.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 74:16:@37549.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 77:19:@37553.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 73:20:@37547.4]
  assign regs_305_clock = clock; // @[:@37556.4]
  assign regs_305_reset = io_reset; // @[:@37557.4 RegFile.scala 75:16:@37564.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 74:16:@37563.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 77:19:@37567.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 73:20:@37561.4]
  assign regs_306_clock = clock; // @[:@37570.4]
  assign regs_306_reset = io_reset; // @[:@37571.4 RegFile.scala 75:16:@37578.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 74:16:@37577.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 77:19:@37581.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 73:20:@37575.4]
  assign regs_307_clock = clock; // @[:@37584.4]
  assign regs_307_reset = io_reset; // @[:@37585.4 RegFile.scala 75:16:@37592.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 74:16:@37591.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 77:19:@37595.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 73:20:@37589.4]
  assign regs_308_clock = clock; // @[:@37598.4]
  assign regs_308_reset = io_reset; // @[:@37599.4 RegFile.scala 75:16:@37606.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 74:16:@37605.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 77:19:@37609.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 73:20:@37603.4]
  assign regs_309_clock = clock; // @[:@37612.4]
  assign regs_309_reset = io_reset; // @[:@37613.4 RegFile.scala 75:16:@37620.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 74:16:@37619.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 77:19:@37623.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 73:20:@37617.4]
  assign regs_310_clock = clock; // @[:@37626.4]
  assign regs_310_reset = io_reset; // @[:@37627.4 RegFile.scala 75:16:@37634.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 74:16:@37633.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 77:19:@37637.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 73:20:@37631.4]
  assign regs_311_clock = clock; // @[:@37640.4]
  assign regs_311_reset = io_reset; // @[:@37641.4 RegFile.scala 75:16:@37648.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 74:16:@37647.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 77:19:@37651.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 73:20:@37645.4]
  assign regs_312_clock = clock; // @[:@37654.4]
  assign regs_312_reset = io_reset; // @[:@37655.4 RegFile.scala 75:16:@37662.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 74:16:@37661.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 77:19:@37665.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 73:20:@37659.4]
  assign regs_313_clock = clock; // @[:@37668.4]
  assign regs_313_reset = io_reset; // @[:@37669.4 RegFile.scala 75:16:@37676.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 74:16:@37675.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 77:19:@37679.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 73:20:@37673.4]
  assign regs_314_clock = clock; // @[:@37682.4]
  assign regs_314_reset = io_reset; // @[:@37683.4 RegFile.scala 75:16:@37690.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 74:16:@37689.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 77:19:@37693.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 73:20:@37687.4]
  assign regs_315_clock = clock; // @[:@37696.4]
  assign regs_315_reset = io_reset; // @[:@37697.4 RegFile.scala 75:16:@37704.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 74:16:@37703.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 77:19:@37707.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 73:20:@37701.4]
  assign regs_316_clock = clock; // @[:@37710.4]
  assign regs_316_reset = io_reset; // @[:@37711.4 RegFile.scala 75:16:@37718.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 74:16:@37717.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 77:19:@37721.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 73:20:@37715.4]
  assign regs_317_clock = clock; // @[:@37724.4]
  assign regs_317_reset = io_reset; // @[:@37725.4 RegFile.scala 75:16:@37732.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 74:16:@37731.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 77:19:@37735.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 73:20:@37729.4]
  assign regs_318_clock = clock; // @[:@37738.4]
  assign regs_318_reset = io_reset; // @[:@37739.4 RegFile.scala 75:16:@37746.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 74:16:@37745.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 77:19:@37749.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 73:20:@37743.4]
  assign regs_319_clock = clock; // @[:@37752.4]
  assign regs_319_reset = io_reset; // @[:@37753.4 RegFile.scala 75:16:@37760.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 74:16:@37759.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 77:19:@37763.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 73:20:@37757.4]
  assign regs_320_clock = clock; // @[:@37766.4]
  assign regs_320_reset = io_reset; // @[:@37767.4 RegFile.scala 75:16:@37774.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 74:16:@37773.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 77:19:@37777.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 73:20:@37771.4]
  assign regs_321_clock = clock; // @[:@37780.4]
  assign regs_321_reset = io_reset; // @[:@37781.4 RegFile.scala 75:16:@37788.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 74:16:@37787.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 77:19:@37791.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 73:20:@37785.4]
  assign regs_322_clock = clock; // @[:@37794.4]
  assign regs_322_reset = io_reset; // @[:@37795.4 RegFile.scala 75:16:@37802.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 74:16:@37801.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 77:19:@37805.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 73:20:@37799.4]
  assign regs_323_clock = clock; // @[:@37808.4]
  assign regs_323_reset = io_reset; // @[:@37809.4 RegFile.scala 75:16:@37816.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 74:16:@37815.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 77:19:@37819.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 73:20:@37813.4]
  assign regs_324_clock = clock; // @[:@37822.4]
  assign regs_324_reset = io_reset; // @[:@37823.4 RegFile.scala 75:16:@37830.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 74:16:@37829.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 77:19:@37833.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 73:20:@37827.4]
  assign regs_325_clock = clock; // @[:@37836.4]
  assign regs_325_reset = io_reset; // @[:@37837.4 RegFile.scala 75:16:@37844.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 74:16:@37843.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 77:19:@37847.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 73:20:@37841.4]
  assign regs_326_clock = clock; // @[:@37850.4]
  assign regs_326_reset = io_reset; // @[:@37851.4 RegFile.scala 75:16:@37858.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 74:16:@37857.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 77:19:@37861.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 73:20:@37855.4]
  assign regs_327_clock = clock; // @[:@37864.4]
  assign regs_327_reset = io_reset; // @[:@37865.4 RegFile.scala 75:16:@37872.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 74:16:@37871.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 77:19:@37875.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 73:20:@37869.4]
  assign regs_328_clock = clock; // @[:@37878.4]
  assign regs_328_reset = io_reset; // @[:@37879.4 RegFile.scala 75:16:@37886.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 74:16:@37885.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 77:19:@37889.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 73:20:@37883.4]
  assign regs_329_clock = clock; // @[:@37892.4]
  assign regs_329_reset = io_reset; // @[:@37893.4 RegFile.scala 75:16:@37900.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 74:16:@37899.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 77:19:@37903.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 73:20:@37897.4]
  assign regs_330_clock = clock; // @[:@37906.4]
  assign regs_330_reset = io_reset; // @[:@37907.4 RegFile.scala 75:16:@37914.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 74:16:@37913.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 77:19:@37917.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 73:20:@37911.4]
  assign regs_331_clock = clock; // @[:@37920.4]
  assign regs_331_reset = io_reset; // @[:@37921.4 RegFile.scala 75:16:@37928.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 74:16:@37927.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 77:19:@37931.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 73:20:@37925.4]
  assign regs_332_clock = clock; // @[:@37934.4]
  assign regs_332_reset = io_reset; // @[:@37935.4 RegFile.scala 75:16:@37942.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 74:16:@37941.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 77:19:@37945.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 73:20:@37939.4]
  assign regs_333_clock = clock; // @[:@37948.4]
  assign regs_333_reset = io_reset; // @[:@37949.4 RegFile.scala 75:16:@37956.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 74:16:@37955.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 77:19:@37959.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 73:20:@37953.4]
  assign regs_334_clock = clock; // @[:@37962.4]
  assign regs_334_reset = io_reset; // @[:@37963.4 RegFile.scala 75:16:@37970.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 74:16:@37969.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 77:19:@37973.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 73:20:@37967.4]
  assign regs_335_clock = clock; // @[:@37976.4]
  assign regs_335_reset = io_reset; // @[:@37977.4 RegFile.scala 75:16:@37984.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 74:16:@37983.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 77:19:@37987.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 73:20:@37981.4]
  assign regs_336_clock = clock; // @[:@37990.4]
  assign regs_336_reset = io_reset; // @[:@37991.4 RegFile.scala 75:16:@37998.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 74:16:@37997.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 77:19:@38001.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 73:20:@37995.4]
  assign regs_337_clock = clock; // @[:@38004.4]
  assign regs_337_reset = io_reset; // @[:@38005.4 RegFile.scala 75:16:@38012.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 74:16:@38011.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 77:19:@38015.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 73:20:@38009.4]
  assign regs_338_clock = clock; // @[:@38018.4]
  assign regs_338_reset = io_reset; // @[:@38019.4 RegFile.scala 75:16:@38026.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 74:16:@38025.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 77:19:@38029.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 73:20:@38023.4]
  assign regs_339_clock = clock; // @[:@38032.4]
  assign regs_339_reset = io_reset; // @[:@38033.4 RegFile.scala 75:16:@38040.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 74:16:@38039.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 77:19:@38043.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 73:20:@38037.4]
  assign regs_340_clock = clock; // @[:@38046.4]
  assign regs_340_reset = io_reset; // @[:@38047.4 RegFile.scala 75:16:@38054.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 74:16:@38053.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 77:19:@38057.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 73:20:@38051.4]
  assign regs_341_clock = clock; // @[:@38060.4]
  assign regs_341_reset = io_reset; // @[:@38061.4 RegFile.scala 75:16:@38068.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 74:16:@38067.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 77:19:@38071.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 73:20:@38065.4]
  assign regs_342_clock = clock; // @[:@38074.4]
  assign regs_342_reset = io_reset; // @[:@38075.4 RegFile.scala 75:16:@38082.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 74:16:@38081.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 77:19:@38085.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 73:20:@38079.4]
  assign regs_343_clock = clock; // @[:@38088.4]
  assign regs_343_reset = io_reset; // @[:@38089.4 RegFile.scala 75:16:@38096.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 74:16:@38095.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 77:19:@38099.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 73:20:@38093.4]
  assign regs_344_clock = clock; // @[:@38102.4]
  assign regs_344_reset = io_reset; // @[:@38103.4 RegFile.scala 75:16:@38110.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 74:16:@38109.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 77:19:@38113.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 73:20:@38107.4]
  assign regs_345_clock = clock; // @[:@38116.4]
  assign regs_345_reset = io_reset; // @[:@38117.4 RegFile.scala 75:16:@38124.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 74:16:@38123.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 77:19:@38127.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 73:20:@38121.4]
  assign regs_346_clock = clock; // @[:@38130.4]
  assign regs_346_reset = io_reset; // @[:@38131.4 RegFile.scala 75:16:@38138.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 74:16:@38137.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 77:19:@38141.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 73:20:@38135.4]
  assign regs_347_clock = clock; // @[:@38144.4]
  assign regs_347_reset = io_reset; // @[:@38145.4 RegFile.scala 75:16:@38152.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 74:16:@38151.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 77:19:@38155.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 73:20:@38149.4]
  assign regs_348_clock = clock; // @[:@38158.4]
  assign regs_348_reset = io_reset; // @[:@38159.4 RegFile.scala 75:16:@38166.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 74:16:@38165.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 77:19:@38169.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 73:20:@38163.4]
  assign regs_349_clock = clock; // @[:@38172.4]
  assign regs_349_reset = io_reset; // @[:@38173.4 RegFile.scala 75:16:@38180.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 74:16:@38179.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 77:19:@38183.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 73:20:@38177.4]
  assign regs_350_clock = clock; // @[:@38186.4]
  assign regs_350_reset = io_reset; // @[:@38187.4 RegFile.scala 75:16:@38194.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 74:16:@38193.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 77:19:@38197.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 73:20:@38191.4]
  assign regs_351_clock = clock; // @[:@38200.4]
  assign regs_351_reset = io_reset; // @[:@38201.4 RegFile.scala 75:16:@38208.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 74:16:@38207.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 77:19:@38211.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 73:20:@38205.4]
  assign regs_352_clock = clock; // @[:@38214.4]
  assign regs_352_reset = io_reset; // @[:@38215.4 RegFile.scala 75:16:@38222.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 74:16:@38221.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 77:19:@38225.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 73:20:@38219.4]
  assign regs_353_clock = clock; // @[:@38228.4]
  assign regs_353_reset = io_reset; // @[:@38229.4 RegFile.scala 75:16:@38236.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 74:16:@38235.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 77:19:@38239.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 73:20:@38233.4]
  assign regs_354_clock = clock; // @[:@38242.4]
  assign regs_354_reset = io_reset; // @[:@38243.4 RegFile.scala 75:16:@38250.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 74:16:@38249.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 77:19:@38253.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 73:20:@38247.4]
  assign regs_355_clock = clock; // @[:@38256.4]
  assign regs_355_reset = io_reset; // @[:@38257.4 RegFile.scala 75:16:@38264.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 74:16:@38263.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 77:19:@38267.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 73:20:@38261.4]
  assign regs_356_clock = clock; // @[:@38270.4]
  assign regs_356_reset = io_reset; // @[:@38271.4 RegFile.scala 75:16:@38278.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 74:16:@38277.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 77:19:@38281.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 73:20:@38275.4]
  assign regs_357_clock = clock; // @[:@38284.4]
  assign regs_357_reset = io_reset; // @[:@38285.4 RegFile.scala 75:16:@38292.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 74:16:@38291.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 77:19:@38295.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 73:20:@38289.4]
  assign regs_358_clock = clock; // @[:@38298.4]
  assign regs_358_reset = io_reset; // @[:@38299.4 RegFile.scala 75:16:@38306.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 74:16:@38305.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 77:19:@38309.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 73:20:@38303.4]
  assign regs_359_clock = clock; // @[:@38312.4]
  assign regs_359_reset = io_reset; // @[:@38313.4 RegFile.scala 75:16:@38320.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 74:16:@38319.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 77:19:@38323.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 73:20:@38317.4]
  assign regs_360_clock = clock; // @[:@38326.4]
  assign regs_360_reset = io_reset; // @[:@38327.4 RegFile.scala 75:16:@38334.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 74:16:@38333.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 77:19:@38337.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 73:20:@38331.4]
  assign regs_361_clock = clock; // @[:@38340.4]
  assign regs_361_reset = io_reset; // @[:@38341.4 RegFile.scala 75:16:@38348.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 74:16:@38347.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 77:19:@38351.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 73:20:@38345.4]
  assign regs_362_clock = clock; // @[:@38354.4]
  assign regs_362_reset = io_reset; // @[:@38355.4 RegFile.scala 75:16:@38362.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 74:16:@38361.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 77:19:@38365.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 73:20:@38359.4]
  assign regs_363_clock = clock; // @[:@38368.4]
  assign regs_363_reset = io_reset; // @[:@38369.4 RegFile.scala 75:16:@38376.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 74:16:@38375.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 77:19:@38379.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 73:20:@38373.4]
  assign regs_364_clock = clock; // @[:@38382.4]
  assign regs_364_reset = io_reset; // @[:@38383.4 RegFile.scala 75:16:@38390.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 74:16:@38389.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 77:19:@38393.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 73:20:@38387.4]
  assign regs_365_clock = clock; // @[:@38396.4]
  assign regs_365_reset = io_reset; // @[:@38397.4 RegFile.scala 75:16:@38404.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 74:16:@38403.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 77:19:@38407.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 73:20:@38401.4]
  assign regs_366_clock = clock; // @[:@38410.4]
  assign regs_366_reset = io_reset; // @[:@38411.4 RegFile.scala 75:16:@38418.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 74:16:@38417.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 77:19:@38421.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 73:20:@38415.4]
  assign regs_367_clock = clock; // @[:@38424.4]
  assign regs_367_reset = io_reset; // @[:@38425.4 RegFile.scala 75:16:@38432.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 74:16:@38431.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 77:19:@38435.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 73:20:@38429.4]
  assign regs_368_clock = clock; // @[:@38438.4]
  assign regs_368_reset = io_reset; // @[:@38439.4 RegFile.scala 75:16:@38446.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 74:16:@38445.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 77:19:@38449.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 73:20:@38443.4]
  assign regs_369_clock = clock; // @[:@38452.4]
  assign regs_369_reset = io_reset; // @[:@38453.4 RegFile.scala 75:16:@38460.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 74:16:@38459.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 77:19:@38463.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 73:20:@38457.4]
  assign regs_370_clock = clock; // @[:@38466.4]
  assign regs_370_reset = io_reset; // @[:@38467.4 RegFile.scala 75:16:@38474.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 74:16:@38473.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 77:19:@38477.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 73:20:@38471.4]
  assign regs_371_clock = clock; // @[:@38480.4]
  assign regs_371_reset = io_reset; // @[:@38481.4 RegFile.scala 75:16:@38488.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 74:16:@38487.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 77:19:@38491.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 73:20:@38485.4]
  assign regs_372_clock = clock; // @[:@38494.4]
  assign regs_372_reset = io_reset; // @[:@38495.4 RegFile.scala 75:16:@38502.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 74:16:@38501.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 77:19:@38505.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 73:20:@38499.4]
  assign regs_373_clock = clock; // @[:@38508.4]
  assign regs_373_reset = io_reset; // @[:@38509.4 RegFile.scala 75:16:@38516.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 74:16:@38515.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 77:19:@38519.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 73:20:@38513.4]
  assign regs_374_clock = clock; // @[:@38522.4]
  assign regs_374_reset = io_reset; // @[:@38523.4 RegFile.scala 75:16:@38530.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 74:16:@38529.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 77:19:@38533.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 73:20:@38527.4]
  assign regs_375_clock = clock; // @[:@38536.4]
  assign regs_375_reset = io_reset; // @[:@38537.4 RegFile.scala 75:16:@38544.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 74:16:@38543.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 77:19:@38547.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 73:20:@38541.4]
  assign regs_376_clock = clock; // @[:@38550.4]
  assign regs_376_reset = io_reset; // @[:@38551.4 RegFile.scala 75:16:@38558.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 74:16:@38557.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 77:19:@38561.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 73:20:@38555.4]
  assign regs_377_clock = clock; // @[:@38564.4]
  assign regs_377_reset = io_reset; // @[:@38565.4 RegFile.scala 75:16:@38572.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 74:16:@38571.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 77:19:@38575.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 73:20:@38569.4]
  assign regs_378_clock = clock; // @[:@38578.4]
  assign regs_378_reset = io_reset; // @[:@38579.4 RegFile.scala 75:16:@38586.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 74:16:@38585.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 77:19:@38589.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 73:20:@38583.4]
  assign regs_379_clock = clock; // @[:@38592.4]
  assign regs_379_reset = io_reset; // @[:@38593.4 RegFile.scala 75:16:@38600.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 74:16:@38599.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 77:19:@38603.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 73:20:@38597.4]
  assign regs_380_clock = clock; // @[:@38606.4]
  assign regs_380_reset = io_reset; // @[:@38607.4 RegFile.scala 75:16:@38614.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 74:16:@38613.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 77:19:@38617.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 73:20:@38611.4]
  assign regs_381_clock = clock; // @[:@38620.4]
  assign regs_381_reset = io_reset; // @[:@38621.4 RegFile.scala 75:16:@38628.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 74:16:@38627.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 77:19:@38631.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 73:20:@38625.4]
  assign regs_382_clock = clock; // @[:@38634.4]
  assign regs_382_reset = io_reset; // @[:@38635.4 RegFile.scala 75:16:@38642.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 74:16:@38641.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 77:19:@38645.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 73:20:@38639.4]
  assign regs_383_clock = clock; // @[:@38648.4]
  assign regs_383_reset = io_reset; // @[:@38649.4 RegFile.scala 75:16:@38656.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 74:16:@38655.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 77:19:@38659.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 73:20:@38653.4]
  assign regs_384_clock = clock; // @[:@38662.4]
  assign regs_384_reset = io_reset; // @[:@38663.4 RegFile.scala 75:16:@38670.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 74:16:@38669.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 77:19:@38673.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 73:20:@38667.4]
  assign regs_385_clock = clock; // @[:@38676.4]
  assign regs_385_reset = io_reset; // @[:@38677.4 RegFile.scala 75:16:@38684.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 74:16:@38683.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 77:19:@38687.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 73:20:@38681.4]
  assign regs_386_clock = clock; // @[:@38690.4]
  assign regs_386_reset = io_reset; // @[:@38691.4 RegFile.scala 75:16:@38698.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 74:16:@38697.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 77:19:@38701.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 73:20:@38695.4]
  assign regs_387_clock = clock; // @[:@38704.4]
  assign regs_387_reset = io_reset; // @[:@38705.4 RegFile.scala 75:16:@38712.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 74:16:@38711.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 77:19:@38715.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 73:20:@38709.4]
  assign regs_388_clock = clock; // @[:@38718.4]
  assign regs_388_reset = io_reset; // @[:@38719.4 RegFile.scala 75:16:@38726.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 74:16:@38725.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 77:19:@38729.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 73:20:@38723.4]
  assign regs_389_clock = clock; // @[:@38732.4]
  assign regs_389_reset = io_reset; // @[:@38733.4 RegFile.scala 75:16:@38740.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 74:16:@38739.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 77:19:@38743.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 73:20:@38737.4]
  assign regs_390_clock = clock; // @[:@38746.4]
  assign regs_390_reset = io_reset; // @[:@38747.4 RegFile.scala 75:16:@38754.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 74:16:@38753.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 77:19:@38757.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 73:20:@38751.4]
  assign regs_391_clock = clock; // @[:@38760.4]
  assign regs_391_reset = io_reset; // @[:@38761.4 RegFile.scala 75:16:@38768.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 74:16:@38767.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 77:19:@38771.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 73:20:@38765.4]
  assign regs_392_clock = clock; // @[:@38774.4]
  assign regs_392_reset = io_reset; // @[:@38775.4 RegFile.scala 75:16:@38782.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 74:16:@38781.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 77:19:@38785.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 73:20:@38779.4]
  assign regs_393_clock = clock; // @[:@38788.4]
  assign regs_393_reset = io_reset; // @[:@38789.4 RegFile.scala 75:16:@38796.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 74:16:@38795.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 77:19:@38799.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 73:20:@38793.4]
  assign regs_394_clock = clock; // @[:@38802.4]
  assign regs_394_reset = io_reset; // @[:@38803.4 RegFile.scala 75:16:@38810.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 74:16:@38809.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 77:19:@38813.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 73:20:@38807.4]
  assign regs_395_clock = clock; // @[:@38816.4]
  assign regs_395_reset = io_reset; // @[:@38817.4 RegFile.scala 75:16:@38824.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 74:16:@38823.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 77:19:@38827.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 73:20:@38821.4]
  assign regs_396_clock = clock; // @[:@38830.4]
  assign regs_396_reset = io_reset; // @[:@38831.4 RegFile.scala 75:16:@38838.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 74:16:@38837.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 77:19:@38841.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 73:20:@38835.4]
  assign regs_397_clock = clock; // @[:@38844.4]
  assign regs_397_reset = io_reset; // @[:@38845.4 RegFile.scala 75:16:@38852.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 74:16:@38851.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 77:19:@38855.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 73:20:@38849.4]
  assign regs_398_clock = clock; // @[:@38858.4]
  assign regs_398_reset = io_reset; // @[:@38859.4 RegFile.scala 75:16:@38866.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 74:16:@38865.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 77:19:@38869.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 73:20:@38863.4]
  assign regs_399_clock = clock; // @[:@38872.4]
  assign regs_399_reset = io_reset; // @[:@38873.4 RegFile.scala 75:16:@38880.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 74:16:@38879.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 77:19:@38883.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 73:20:@38877.4]
  assign regs_400_clock = clock; // @[:@38886.4]
  assign regs_400_reset = io_reset; // @[:@38887.4 RegFile.scala 75:16:@38894.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 74:16:@38893.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 77:19:@38897.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 73:20:@38891.4]
  assign regs_401_clock = clock; // @[:@38900.4]
  assign regs_401_reset = io_reset; // @[:@38901.4 RegFile.scala 75:16:@38908.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 74:16:@38907.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 77:19:@38911.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 73:20:@38905.4]
  assign regs_402_clock = clock; // @[:@38914.4]
  assign regs_402_reset = io_reset; // @[:@38915.4 RegFile.scala 75:16:@38922.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 74:16:@38921.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 77:19:@38925.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 73:20:@38919.4]
  assign regs_403_clock = clock; // @[:@38928.4]
  assign regs_403_reset = io_reset; // @[:@38929.4 RegFile.scala 75:16:@38936.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 74:16:@38935.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 77:19:@38939.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 73:20:@38933.4]
  assign regs_404_clock = clock; // @[:@38942.4]
  assign regs_404_reset = io_reset; // @[:@38943.4 RegFile.scala 75:16:@38950.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 74:16:@38949.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 77:19:@38953.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 73:20:@38947.4]
  assign regs_405_clock = clock; // @[:@38956.4]
  assign regs_405_reset = io_reset; // @[:@38957.4 RegFile.scala 75:16:@38964.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 74:16:@38963.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 77:19:@38967.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 73:20:@38961.4]
  assign regs_406_clock = clock; // @[:@38970.4]
  assign regs_406_reset = io_reset; // @[:@38971.4 RegFile.scala 75:16:@38978.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 74:16:@38977.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 77:19:@38981.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 73:20:@38975.4]
  assign regs_407_clock = clock; // @[:@38984.4]
  assign regs_407_reset = io_reset; // @[:@38985.4 RegFile.scala 75:16:@38992.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 74:16:@38991.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 77:19:@38995.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 73:20:@38989.4]
  assign regs_408_clock = clock; // @[:@38998.4]
  assign regs_408_reset = io_reset; // @[:@38999.4 RegFile.scala 75:16:@39006.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 74:16:@39005.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 77:19:@39009.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 73:20:@39003.4]
  assign regs_409_clock = clock; // @[:@39012.4]
  assign regs_409_reset = io_reset; // @[:@39013.4 RegFile.scala 75:16:@39020.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 74:16:@39019.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 77:19:@39023.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 73:20:@39017.4]
  assign regs_410_clock = clock; // @[:@39026.4]
  assign regs_410_reset = io_reset; // @[:@39027.4 RegFile.scala 75:16:@39034.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 74:16:@39033.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 77:19:@39037.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 73:20:@39031.4]
  assign regs_411_clock = clock; // @[:@39040.4]
  assign regs_411_reset = io_reset; // @[:@39041.4 RegFile.scala 75:16:@39048.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 74:16:@39047.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 77:19:@39051.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 73:20:@39045.4]
  assign regs_412_clock = clock; // @[:@39054.4]
  assign regs_412_reset = io_reset; // @[:@39055.4 RegFile.scala 75:16:@39062.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 74:16:@39061.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 77:19:@39065.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 73:20:@39059.4]
  assign regs_413_clock = clock; // @[:@39068.4]
  assign regs_413_reset = io_reset; // @[:@39069.4 RegFile.scala 75:16:@39076.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 74:16:@39075.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 77:19:@39079.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 73:20:@39073.4]
  assign regs_414_clock = clock; // @[:@39082.4]
  assign regs_414_reset = io_reset; // @[:@39083.4 RegFile.scala 75:16:@39090.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 74:16:@39089.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 77:19:@39093.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 73:20:@39087.4]
  assign regs_415_clock = clock; // @[:@39096.4]
  assign regs_415_reset = io_reset; // @[:@39097.4 RegFile.scala 75:16:@39104.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 74:16:@39103.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 77:19:@39107.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 73:20:@39101.4]
  assign regs_416_clock = clock; // @[:@39110.4]
  assign regs_416_reset = io_reset; // @[:@39111.4 RegFile.scala 75:16:@39118.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 74:16:@39117.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 77:19:@39121.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 73:20:@39115.4]
  assign regs_417_clock = clock; // @[:@39124.4]
  assign regs_417_reset = io_reset; // @[:@39125.4 RegFile.scala 75:16:@39132.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 74:16:@39131.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 77:19:@39135.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 73:20:@39129.4]
  assign regs_418_clock = clock; // @[:@39138.4]
  assign regs_418_reset = io_reset; // @[:@39139.4 RegFile.scala 75:16:@39146.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 74:16:@39145.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 77:19:@39149.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 73:20:@39143.4]
  assign regs_419_clock = clock; // @[:@39152.4]
  assign regs_419_reset = io_reset; // @[:@39153.4 RegFile.scala 75:16:@39160.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 74:16:@39159.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 77:19:@39163.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 73:20:@39157.4]
  assign regs_420_clock = clock; // @[:@39166.4]
  assign regs_420_reset = io_reset; // @[:@39167.4 RegFile.scala 75:16:@39174.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 74:16:@39173.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 77:19:@39177.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 73:20:@39171.4]
  assign regs_421_clock = clock; // @[:@39180.4]
  assign regs_421_reset = io_reset; // @[:@39181.4 RegFile.scala 75:16:@39188.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 74:16:@39187.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 77:19:@39191.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 73:20:@39185.4]
  assign regs_422_clock = clock; // @[:@39194.4]
  assign regs_422_reset = io_reset; // @[:@39195.4 RegFile.scala 75:16:@39202.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 74:16:@39201.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 77:19:@39205.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 73:20:@39199.4]
  assign regs_423_clock = clock; // @[:@39208.4]
  assign regs_423_reset = io_reset; // @[:@39209.4 RegFile.scala 75:16:@39216.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 74:16:@39215.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 77:19:@39219.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 73:20:@39213.4]
  assign regs_424_clock = clock; // @[:@39222.4]
  assign regs_424_reset = io_reset; // @[:@39223.4 RegFile.scala 75:16:@39230.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 74:16:@39229.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 77:19:@39233.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 73:20:@39227.4]
  assign regs_425_clock = clock; // @[:@39236.4]
  assign regs_425_reset = io_reset; // @[:@39237.4 RegFile.scala 75:16:@39244.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 74:16:@39243.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 77:19:@39247.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 73:20:@39241.4]
  assign regs_426_clock = clock; // @[:@39250.4]
  assign regs_426_reset = io_reset; // @[:@39251.4 RegFile.scala 75:16:@39258.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 74:16:@39257.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 77:19:@39261.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 73:20:@39255.4]
  assign regs_427_clock = clock; // @[:@39264.4]
  assign regs_427_reset = io_reset; // @[:@39265.4 RegFile.scala 75:16:@39272.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 74:16:@39271.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 77:19:@39275.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 73:20:@39269.4]
  assign regs_428_clock = clock; // @[:@39278.4]
  assign regs_428_reset = io_reset; // @[:@39279.4 RegFile.scala 75:16:@39286.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 74:16:@39285.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 77:19:@39289.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 73:20:@39283.4]
  assign regs_429_clock = clock; // @[:@39292.4]
  assign regs_429_reset = io_reset; // @[:@39293.4 RegFile.scala 75:16:@39300.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 74:16:@39299.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 77:19:@39303.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 73:20:@39297.4]
  assign regs_430_clock = clock; // @[:@39306.4]
  assign regs_430_reset = io_reset; // @[:@39307.4 RegFile.scala 75:16:@39314.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 74:16:@39313.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 77:19:@39317.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 73:20:@39311.4]
  assign regs_431_clock = clock; // @[:@39320.4]
  assign regs_431_reset = io_reset; // @[:@39321.4 RegFile.scala 75:16:@39328.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 74:16:@39327.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 77:19:@39331.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 73:20:@39325.4]
  assign regs_432_clock = clock; // @[:@39334.4]
  assign regs_432_reset = io_reset; // @[:@39335.4 RegFile.scala 75:16:@39342.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 74:16:@39341.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 77:19:@39345.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 73:20:@39339.4]
  assign regs_433_clock = clock; // @[:@39348.4]
  assign regs_433_reset = io_reset; // @[:@39349.4 RegFile.scala 75:16:@39356.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 74:16:@39355.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 77:19:@39359.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 73:20:@39353.4]
  assign regs_434_clock = clock; // @[:@39362.4]
  assign regs_434_reset = io_reset; // @[:@39363.4 RegFile.scala 75:16:@39370.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 74:16:@39369.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 77:19:@39373.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 73:20:@39367.4]
  assign regs_435_clock = clock; // @[:@39376.4]
  assign regs_435_reset = io_reset; // @[:@39377.4 RegFile.scala 75:16:@39384.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 74:16:@39383.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 77:19:@39387.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 73:20:@39381.4]
  assign regs_436_clock = clock; // @[:@39390.4]
  assign regs_436_reset = io_reset; // @[:@39391.4 RegFile.scala 75:16:@39398.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 74:16:@39397.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 77:19:@39401.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 73:20:@39395.4]
  assign regs_437_clock = clock; // @[:@39404.4]
  assign regs_437_reset = io_reset; // @[:@39405.4 RegFile.scala 75:16:@39412.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 74:16:@39411.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 77:19:@39415.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 73:20:@39409.4]
  assign regs_438_clock = clock; // @[:@39418.4]
  assign regs_438_reset = io_reset; // @[:@39419.4 RegFile.scala 75:16:@39426.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 74:16:@39425.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 77:19:@39429.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 73:20:@39423.4]
  assign regs_439_clock = clock; // @[:@39432.4]
  assign regs_439_reset = io_reset; // @[:@39433.4 RegFile.scala 75:16:@39440.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 74:16:@39439.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 77:19:@39443.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 73:20:@39437.4]
  assign regs_440_clock = clock; // @[:@39446.4]
  assign regs_440_reset = io_reset; // @[:@39447.4 RegFile.scala 75:16:@39454.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 74:16:@39453.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 77:19:@39457.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 73:20:@39451.4]
  assign regs_441_clock = clock; // @[:@39460.4]
  assign regs_441_reset = io_reset; // @[:@39461.4 RegFile.scala 75:16:@39468.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 74:16:@39467.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 77:19:@39471.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 73:20:@39465.4]
  assign regs_442_clock = clock; // @[:@39474.4]
  assign regs_442_reset = io_reset; // @[:@39475.4 RegFile.scala 75:16:@39482.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 74:16:@39481.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 77:19:@39485.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 73:20:@39479.4]
  assign regs_443_clock = clock; // @[:@39488.4]
  assign regs_443_reset = io_reset; // @[:@39489.4 RegFile.scala 75:16:@39496.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 74:16:@39495.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 77:19:@39499.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 73:20:@39493.4]
  assign regs_444_clock = clock; // @[:@39502.4]
  assign regs_444_reset = io_reset; // @[:@39503.4 RegFile.scala 75:16:@39510.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 74:16:@39509.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 77:19:@39513.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 73:20:@39507.4]
  assign regs_445_clock = clock; // @[:@39516.4]
  assign regs_445_reset = io_reset; // @[:@39517.4 RegFile.scala 75:16:@39524.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 74:16:@39523.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 77:19:@39527.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 73:20:@39521.4]
  assign regs_446_clock = clock; // @[:@39530.4]
  assign regs_446_reset = io_reset; // @[:@39531.4 RegFile.scala 75:16:@39538.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 74:16:@39537.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 77:19:@39541.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 73:20:@39535.4]
  assign regs_447_clock = clock; // @[:@39544.4]
  assign regs_447_reset = io_reset; // @[:@39545.4 RegFile.scala 75:16:@39552.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 74:16:@39551.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 77:19:@39555.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 73:20:@39549.4]
  assign regs_448_clock = clock; // @[:@39558.4]
  assign regs_448_reset = io_reset; // @[:@39559.4 RegFile.scala 75:16:@39566.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 74:16:@39565.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 77:19:@39569.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 73:20:@39563.4]
  assign regs_449_clock = clock; // @[:@39572.4]
  assign regs_449_reset = io_reset; // @[:@39573.4 RegFile.scala 75:16:@39580.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 74:16:@39579.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 77:19:@39583.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 73:20:@39577.4]
  assign regs_450_clock = clock; // @[:@39586.4]
  assign regs_450_reset = io_reset; // @[:@39587.4 RegFile.scala 75:16:@39594.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 74:16:@39593.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 77:19:@39597.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 73:20:@39591.4]
  assign regs_451_clock = clock; // @[:@39600.4]
  assign regs_451_reset = io_reset; // @[:@39601.4 RegFile.scala 75:16:@39608.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 74:16:@39607.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 77:19:@39611.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 73:20:@39605.4]
  assign regs_452_clock = clock; // @[:@39614.4]
  assign regs_452_reset = io_reset; // @[:@39615.4 RegFile.scala 75:16:@39622.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 74:16:@39621.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 77:19:@39625.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 73:20:@39619.4]
  assign regs_453_clock = clock; // @[:@39628.4]
  assign regs_453_reset = io_reset; // @[:@39629.4 RegFile.scala 75:16:@39636.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 74:16:@39635.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 77:19:@39639.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 73:20:@39633.4]
  assign regs_454_clock = clock; // @[:@39642.4]
  assign regs_454_reset = io_reset; // @[:@39643.4 RegFile.scala 75:16:@39650.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 74:16:@39649.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 77:19:@39653.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 73:20:@39647.4]
  assign regs_455_clock = clock; // @[:@39656.4]
  assign regs_455_reset = io_reset; // @[:@39657.4 RegFile.scala 75:16:@39664.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 74:16:@39663.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 77:19:@39667.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 73:20:@39661.4]
  assign regs_456_clock = clock; // @[:@39670.4]
  assign regs_456_reset = io_reset; // @[:@39671.4 RegFile.scala 75:16:@39678.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 74:16:@39677.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 77:19:@39681.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 73:20:@39675.4]
  assign regs_457_clock = clock; // @[:@39684.4]
  assign regs_457_reset = io_reset; // @[:@39685.4 RegFile.scala 75:16:@39692.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 74:16:@39691.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 77:19:@39695.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 73:20:@39689.4]
  assign regs_458_clock = clock; // @[:@39698.4]
  assign regs_458_reset = io_reset; // @[:@39699.4 RegFile.scala 75:16:@39706.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 74:16:@39705.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 77:19:@39709.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 73:20:@39703.4]
  assign regs_459_clock = clock; // @[:@39712.4]
  assign regs_459_reset = io_reset; // @[:@39713.4 RegFile.scala 75:16:@39720.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 74:16:@39719.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 77:19:@39723.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 73:20:@39717.4]
  assign regs_460_clock = clock; // @[:@39726.4]
  assign regs_460_reset = io_reset; // @[:@39727.4 RegFile.scala 75:16:@39734.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 74:16:@39733.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 77:19:@39737.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 73:20:@39731.4]
  assign regs_461_clock = clock; // @[:@39740.4]
  assign regs_461_reset = io_reset; // @[:@39741.4 RegFile.scala 75:16:@39748.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 74:16:@39747.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 77:19:@39751.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 73:20:@39745.4]
  assign regs_462_clock = clock; // @[:@39754.4]
  assign regs_462_reset = io_reset; // @[:@39755.4 RegFile.scala 75:16:@39762.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 74:16:@39761.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 77:19:@39765.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 73:20:@39759.4]
  assign regs_463_clock = clock; // @[:@39768.4]
  assign regs_463_reset = io_reset; // @[:@39769.4 RegFile.scala 75:16:@39776.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 74:16:@39775.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 77:19:@39779.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 73:20:@39773.4]
  assign regs_464_clock = clock; // @[:@39782.4]
  assign regs_464_reset = io_reset; // @[:@39783.4 RegFile.scala 75:16:@39790.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 74:16:@39789.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 77:19:@39793.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 73:20:@39787.4]
  assign regs_465_clock = clock; // @[:@39796.4]
  assign regs_465_reset = io_reset; // @[:@39797.4 RegFile.scala 75:16:@39804.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 74:16:@39803.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 77:19:@39807.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 73:20:@39801.4]
  assign regs_466_clock = clock; // @[:@39810.4]
  assign regs_466_reset = io_reset; // @[:@39811.4 RegFile.scala 75:16:@39818.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 74:16:@39817.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 77:19:@39821.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 73:20:@39815.4]
  assign regs_467_clock = clock; // @[:@39824.4]
  assign regs_467_reset = io_reset; // @[:@39825.4 RegFile.scala 75:16:@39832.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 74:16:@39831.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 77:19:@39835.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 73:20:@39829.4]
  assign regs_468_clock = clock; // @[:@39838.4]
  assign regs_468_reset = io_reset; // @[:@39839.4 RegFile.scala 75:16:@39846.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 74:16:@39845.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 77:19:@39849.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 73:20:@39843.4]
  assign regs_469_clock = clock; // @[:@39852.4]
  assign regs_469_reset = io_reset; // @[:@39853.4 RegFile.scala 75:16:@39860.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 74:16:@39859.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 77:19:@39863.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 73:20:@39857.4]
  assign regs_470_clock = clock; // @[:@39866.4]
  assign regs_470_reset = io_reset; // @[:@39867.4 RegFile.scala 75:16:@39874.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 74:16:@39873.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 77:19:@39877.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 73:20:@39871.4]
  assign regs_471_clock = clock; // @[:@39880.4]
  assign regs_471_reset = io_reset; // @[:@39881.4 RegFile.scala 75:16:@39888.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 74:16:@39887.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 77:19:@39891.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 73:20:@39885.4]
  assign regs_472_clock = clock; // @[:@39894.4]
  assign regs_472_reset = io_reset; // @[:@39895.4 RegFile.scala 75:16:@39902.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 74:16:@39901.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 77:19:@39905.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 73:20:@39899.4]
  assign regs_473_clock = clock; // @[:@39908.4]
  assign regs_473_reset = io_reset; // @[:@39909.4 RegFile.scala 75:16:@39916.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 74:16:@39915.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 77:19:@39919.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 73:20:@39913.4]
  assign regs_474_clock = clock; // @[:@39922.4]
  assign regs_474_reset = io_reset; // @[:@39923.4 RegFile.scala 75:16:@39930.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 74:16:@39929.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 77:19:@39933.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 73:20:@39927.4]
  assign regs_475_clock = clock; // @[:@39936.4]
  assign regs_475_reset = io_reset; // @[:@39937.4 RegFile.scala 75:16:@39944.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 74:16:@39943.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 77:19:@39947.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 73:20:@39941.4]
  assign regs_476_clock = clock; // @[:@39950.4]
  assign regs_476_reset = io_reset; // @[:@39951.4 RegFile.scala 75:16:@39958.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 74:16:@39957.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 77:19:@39961.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 73:20:@39955.4]
  assign regs_477_clock = clock; // @[:@39964.4]
  assign regs_477_reset = io_reset; // @[:@39965.4 RegFile.scala 75:16:@39972.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 74:16:@39971.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 77:19:@39975.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 73:20:@39969.4]
  assign regs_478_clock = clock; // @[:@39978.4]
  assign regs_478_reset = io_reset; // @[:@39979.4 RegFile.scala 75:16:@39986.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 74:16:@39985.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 77:19:@39989.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 73:20:@39983.4]
  assign regs_479_clock = clock; // @[:@39992.4]
  assign regs_479_reset = io_reset; // @[:@39993.4 RegFile.scala 75:16:@40000.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 74:16:@39999.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 77:19:@40003.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 73:20:@39997.4]
  assign regs_480_clock = clock; // @[:@40006.4]
  assign regs_480_reset = io_reset; // @[:@40007.4 RegFile.scala 75:16:@40014.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 74:16:@40013.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 77:19:@40017.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 73:20:@40011.4]
  assign regs_481_clock = clock; // @[:@40020.4]
  assign regs_481_reset = io_reset; // @[:@40021.4 RegFile.scala 75:16:@40028.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 74:16:@40027.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 77:19:@40031.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 73:20:@40025.4]
  assign regs_482_clock = clock; // @[:@40034.4]
  assign regs_482_reset = io_reset; // @[:@40035.4 RegFile.scala 75:16:@40042.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 74:16:@40041.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 77:19:@40045.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 73:20:@40039.4]
  assign regs_483_clock = clock; // @[:@40048.4]
  assign regs_483_reset = io_reset; // @[:@40049.4 RegFile.scala 75:16:@40056.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 74:16:@40055.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 77:19:@40059.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 73:20:@40053.4]
  assign regs_484_clock = clock; // @[:@40062.4]
  assign regs_484_reset = io_reset; // @[:@40063.4 RegFile.scala 75:16:@40070.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 74:16:@40069.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 77:19:@40073.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 73:20:@40067.4]
  assign regs_485_clock = clock; // @[:@40076.4]
  assign regs_485_reset = io_reset; // @[:@40077.4 RegFile.scala 75:16:@40084.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 74:16:@40083.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 77:19:@40087.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 73:20:@40081.4]
  assign regs_486_clock = clock; // @[:@40090.4]
  assign regs_486_reset = io_reset; // @[:@40091.4 RegFile.scala 75:16:@40098.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 74:16:@40097.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 77:19:@40101.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 73:20:@40095.4]
  assign regs_487_clock = clock; // @[:@40104.4]
  assign regs_487_reset = io_reset; // @[:@40105.4 RegFile.scala 75:16:@40112.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 74:16:@40111.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 77:19:@40115.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 73:20:@40109.4]
  assign regs_488_clock = clock; // @[:@40118.4]
  assign regs_488_reset = io_reset; // @[:@40119.4 RegFile.scala 75:16:@40126.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 74:16:@40125.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 77:19:@40129.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 73:20:@40123.4]
  assign regs_489_clock = clock; // @[:@40132.4]
  assign regs_489_reset = io_reset; // @[:@40133.4 RegFile.scala 75:16:@40140.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 74:16:@40139.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 77:19:@40143.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 73:20:@40137.4]
  assign regs_490_clock = clock; // @[:@40146.4]
  assign regs_490_reset = io_reset; // @[:@40147.4 RegFile.scala 75:16:@40154.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 74:16:@40153.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 77:19:@40157.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 73:20:@40151.4]
  assign regs_491_clock = clock; // @[:@40160.4]
  assign regs_491_reset = io_reset; // @[:@40161.4 RegFile.scala 75:16:@40168.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 74:16:@40167.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 77:19:@40171.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 73:20:@40165.4]
  assign regs_492_clock = clock; // @[:@40174.4]
  assign regs_492_reset = io_reset; // @[:@40175.4 RegFile.scala 75:16:@40182.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 74:16:@40181.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 77:19:@40185.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 73:20:@40179.4]
  assign regs_493_clock = clock; // @[:@40188.4]
  assign regs_493_reset = io_reset; // @[:@40189.4 RegFile.scala 75:16:@40196.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 74:16:@40195.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 77:19:@40199.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 73:20:@40193.4]
  assign regs_494_clock = clock; // @[:@40202.4]
  assign regs_494_reset = io_reset; // @[:@40203.4 RegFile.scala 75:16:@40210.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 74:16:@40209.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 77:19:@40213.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 73:20:@40207.4]
  assign regs_495_clock = clock; // @[:@40216.4]
  assign regs_495_reset = io_reset; // @[:@40217.4 RegFile.scala 75:16:@40224.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 74:16:@40223.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 77:19:@40227.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 73:20:@40221.4]
  assign regs_496_clock = clock; // @[:@40230.4]
  assign regs_496_reset = io_reset; // @[:@40231.4 RegFile.scala 75:16:@40238.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 74:16:@40237.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 77:19:@40241.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 73:20:@40235.4]
  assign regs_497_clock = clock; // @[:@40244.4]
  assign regs_497_reset = io_reset; // @[:@40245.4 RegFile.scala 75:16:@40252.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 74:16:@40251.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 77:19:@40255.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 73:20:@40249.4]
  assign regs_498_clock = clock; // @[:@40258.4]
  assign regs_498_reset = io_reset; // @[:@40259.4 RegFile.scala 75:16:@40266.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 74:16:@40265.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 77:19:@40269.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 73:20:@40263.4]
  assign regs_499_clock = clock; // @[:@40272.4]
  assign regs_499_reset = io_reset; // @[:@40273.4 RegFile.scala 75:16:@40280.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 74:16:@40279.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 77:19:@40283.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 73:20:@40277.4]
  assign regs_500_clock = clock; // @[:@40286.4]
  assign regs_500_reset = io_reset; // @[:@40287.4 RegFile.scala 75:16:@40294.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 74:16:@40293.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 77:19:@40297.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 73:20:@40291.4]
  assign regs_501_clock = clock; // @[:@40300.4]
  assign regs_501_reset = io_reset; // @[:@40301.4 RegFile.scala 75:16:@40308.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 74:16:@40307.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 77:19:@40311.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 73:20:@40305.4]
  assign regs_502_clock = clock; // @[:@40314.4]
  assign regs_502_reset = io_reset; // @[:@40315.4 RegFile.scala 75:16:@40322.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 74:16:@40321.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 77:19:@40325.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 73:20:@40319.4]
endmodule
module RetimeWrapper_507( // @[:@41359.2]
  input         clock, // @[:@41360.4]
  input         reset, // @[:@41361.4]
  input  [39:0] io_in, // @[:@41362.4]
  output [39:0] io_out // @[:@41362.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@41364.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@41364.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@41377.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@41376.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@41375.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@41374.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@41373.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@41371.4]
endmodule
module FringeFF_503( // @[:@41379.2]
  input         clock, // @[:@41380.4]
  input         reset, // @[:@41381.4]
  input  [39:0] io_in, // @[:@41382.4]
  output [39:0] io_out, // @[:@41382.4]
  input         io_enable // @[:@41382.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 98:22:@41385.4]
  wire  RetimeWrapper_reset; // @[package.scala 98:22:@41385.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 98:22:@41385.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 98:22:@41385.4]
  wire [39:0] _T_18; // @[package.scala 101:25:@41390.4 package.scala 101:25:@41391.4]
  RetimeWrapper_507 RetimeWrapper ( // @[package.scala 98:22:@41385.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 101:25:@41390.4 package.scala 101:25:@41391.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@41402.4]
  assign RetimeWrapper_clock = clock; // @[:@41386.4]
  assign RetimeWrapper_reset = reset; // @[:@41387.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 99:16:@41388.4]
endmodule
module FringeCounter( // @[:@41404.2]
  input   clock, // @[:@41405.4]
  input   reset, // @[:@41406.4]
  input   io_enable, // @[:@41407.4]
  output  io_done // @[:@41407.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@41409.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@41409.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@41409.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@41409.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@41409.4]
  wire [40:0] count; // @[Cat.scala 30:58:@41416.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@41417.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@41418.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@41419.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@41421.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@41409.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@41416.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@41417.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@41418.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@41419.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@41421.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@41432.4]
  assign reg$_clock = clock; // @[:@41410.4]
  assign reg$_reset = reset; // @[:@41411.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@41423.6 FringeCounter.scala 37:15:@41426.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@41414.4]
endmodule
module FringeFF_504( // @[:@41466.2]
  input   clock, // @[:@41467.4]
  input   reset, // @[:@41468.4]
  input   io_in, // @[:@41469.4]
  input   io_reset, // @[:@41469.4]
  output  io_out, // @[:@41469.4]
  input   io_enable // @[:@41469.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 98:22:@41472.4]
  wire  RetimeWrapper_reset; // @[package.scala 98:22:@41472.4]
  wire  RetimeWrapper_io_in; // @[package.scala 98:22:@41472.4]
  wire  RetimeWrapper_io_out; // @[package.scala 98:22:@41472.4]
  wire  _T_18; // @[package.scala 101:25:@41477.4 package.scala 101:25:@41478.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@41483.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 98:22:@41472.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 101:25:@41477.4 package.scala 101:25:@41478.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@41483.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@41489.4]
  assign RetimeWrapper_clock = clock; // @[:@41473.4]
  assign RetimeWrapper_reset = reset; // @[:@41474.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 99:16:@41475.4]
endmodule
module Depulser( // @[:@41491.2]
  input   clock, // @[:@41492.4]
  input   reset, // @[:@41493.4]
  input   io_in, // @[:@41494.4]
  input   io_rst, // @[:@41494.4]
  output  io_out // @[:@41494.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@41496.4]
  wire  r_reset; // @[Depulser.scala 14:17:@41496.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@41496.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@41496.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@41496.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@41496.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@41496.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@41505.4]
  assign r_clock = clock; // @[:@41497.4]
  assign r_reset = reset; // @[:@41498.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@41500.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@41504.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@41503.4]
endmodule
module Fringe( // @[:@41507.2]
  input         clock, // @[:@41508.4]
  input         reset, // @[:@41509.4]
  output        io_enable, // @[:@41510.4]
  input         io_done, // @[:@41510.4]
  output        io_reset, // @[:@41510.4]
  output [63:0] io_argIns_0, // @[:@41510.4]
  input         io_argOuts_0_valid, // @[:@41510.4]
  input  [63:0] io_argOuts_0_bits // @[:@41510.4]
);
  wire  regs_clock; // @[Fringe.scala 116:20:@43315.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@43315.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@43315.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@43315.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@43315.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@43315.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@43315.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@43315.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@43315.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@43315.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@45364.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@45364.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@45364.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@45364.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@45382.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@45382.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@45382.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@45382.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@45382.4]
  wire [63:0] _T_874; // @[:@45341.4 :@45342.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@45343.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@45345.4]
  wire  _T_879; // @[Fringe.scala 134:28:@45351.4]
  wire  _T_883; // @[Fringe.scala 134:42:@45353.4]
  wire  _T_884; // @[Fringe.scala 135:27:@45355.4]
  wire [63:0] _T_894; // @[Fringe.scala 156:22:@45390.4]
  wire  _T_906; // @[Fringe.scala 160:55:@45400.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@45401.4]
  wire  _T_909; // @[Fringe.scala 161:58:@45404.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@45405.4]
  wire [1:0] _T_918; // @[Fringe.scala 171:37:@45413.4]
  RegFile regs ( // @[Fringe.scala 116:20:@43315.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@45364.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@45382.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_874 = regs_io_argIns_1; // @[:@45341.4 :@45342.4]
  assign curStatus_done = _T_874[0]; // @[Fringe.scala 133:45:@45343.4]
  assign curStatus_timeout = _T_874[1]; // @[Fringe.scala 133:45:@45345.4]
  assign _T_879 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@45351.4]
  assign _T_883 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@45353.4]
  assign _T_884 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@45355.4]
  assign _T_894 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@45390.4]
  assign _T_906 = _T_879 & depulser_io_out; // @[Fringe.scala 160:55:@45400.4]
  assign status_bits_done = depulser_io_out ? _T_906 : curStatus_done; // @[Fringe.scala 160:26:@45401.4]
  assign _T_909 = _T_879 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@45404.4]
  assign status_bits_timeout = depulser_io_out ? _T_909 : curStatus_timeout; // @[Fringe.scala 161:29:@45405.4]
  assign _T_918 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@45413.4]
  assign io_enable = _T_879 & _T_883; // @[Fringe.scala 136:13:@45359.4]
  assign io_reset = _T_884 | reset; // @[Fringe.scala 137:12:@45360.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@45381.4]
  assign regs_clock = clock; // @[:@43316.4]
  assign regs_reset = reset; // @[:@43317.4 Fringe.scala 139:14:@45363.4]
  assign regs_io_reset = _T_884 | reset; // @[Fringe.scala 138:17:@45361.4]
  assign regs_io_argOuts_0_valid = depulser_io_out; // @[Fringe.scala 170:23:@45412.4]
  assign regs_io_argOuts_0_bits = {62'h0,_T_918}; // @[Fringe.scala 171:22:@45416.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@45419.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@45418.4]
  assign timeoutCtr_clock = clock; // @[:@45365.4]
  assign timeoutCtr_reset = reset; // @[:@45366.4]
  assign timeoutCtr_io_enable = _T_879 & _T_883; // @[Fringe.scala 149:24:@45380.4]
  assign depulser_clock = clock; // @[:@45383.4]
  assign depulser_reset = reset; // @[:@45384.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@45389.4]
  assign depulser_io_rst = _T_894[0]; // @[Fringe.scala 156:19:@45391.4]
endmodule
module MAGToAXI4Bridge( // @[:@46793.2]
  output [7:0] io_M_AXI_AWLEN, // @[:@46796.4]
  output [7:0] io_M_AXI_ARLEN // @[:@46796.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@46937.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@46938.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@46939.4]
  assign _T_218 = 32'h0 - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@46937.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@46938.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@46939.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@46957.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@46940.4]
endmodule
module FringeZynq( // @[:@47353.2]
  input         clock, // @[:@47354.4]
  input         reset, // @[:@47355.4]
  output [7:0]  io_M_AXI_0_AWLEN, // @[:@47356.4]
  output [7:0]  io_M_AXI_0_ARLEN, // @[:@47356.4]
  output [7:0]  io_M_AXI_1_AWLEN, // @[:@47356.4]
  output [7:0]  io_M_AXI_1_ARLEN, // @[:@47356.4]
  output        io_enable, // @[:@47356.4]
  input         io_done, // @[:@47356.4]
  output        io_reset, // @[:@47356.4]
  output [63:0] io_argIns_0, // @[:@47356.4]
  input         io_argOuts_0_valid, // @[:@47356.4]
  input  [63:0] io_argOuts_0_bits // @[:@47356.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 68:28:@47711.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 68:28:@47711.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 68:28:@47711.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 68:28:@47711.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 68:28:@47711.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 68:28:@47711.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 68:28:@47711.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 68:28:@47711.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 119:27:@48416.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 119:27:@48416.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 119:27:@48556.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 119:27:@48556.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 68:28:@47711.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 119:27:@48416.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 119:27:@48556.4]
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN)
  );
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 121:10:@48552.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 121:10:@48540.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 121:10:@48692.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 121:10:@48680.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 103:13:@48328.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 107:12:@48332.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 109:13:@48333.4]
  assign fringeCommon_clock = clock; // @[:@47712.4]
  assign fringeCommon_reset = reset; // @[:@47713.4 FringeZynq.scala 105:22:@48331.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 104:24:@48329.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 110:27:@48335.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 110:27:@48334.4]
endmodule
module Top( // @[:@48697.2]
  input          clock, // @[:@48698.4]
  input          reset, // @[:@48699.4]
  input          io_raddr, // @[:@48700.4]
  input          io_wen, // @[:@48700.4]
  input          io_waddr, // @[:@48700.4]
  input          io_wdata, // @[:@48700.4]
  output         io_rdata, // @[:@48700.4]
  input  [39:0]  io_S_AXI_AWADDR, // @[:@48700.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@48700.4]
  input          io_S_AXI_AWVALID, // @[:@48700.4]
  output         io_S_AXI_AWREADY, // @[:@48700.4]
  input  [39:0]  io_S_AXI_ARADDR, // @[:@48700.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@48700.4]
  input          io_S_AXI_ARVALID, // @[:@48700.4]
  output         io_S_AXI_ARREADY, // @[:@48700.4]
  input  [63:0]  io_S_AXI_WDATA, // @[:@48700.4]
  input  [7:0]   io_S_AXI_WSTRB, // @[:@48700.4]
  input          io_S_AXI_WVALID, // @[:@48700.4]
  output         io_S_AXI_WREADY, // @[:@48700.4]
  output [63:0]  io_S_AXI_RDATA, // @[:@48700.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@48700.4]
  output         io_S_AXI_RVALID, // @[:@48700.4]
  input          io_S_AXI_RREADY, // @[:@48700.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@48700.4]
  output         io_S_AXI_BVALID, // @[:@48700.4]
  input          io_S_AXI_BREADY, // @[:@48700.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@48700.4]
  output [39:0]  io_M_AXI_0_AWUSER, // @[:@48700.4]
  output [39:0]  io_M_AXI_0_AWADDR, // @[:@48700.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@48700.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@48700.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@48700.4]
  output         io_M_AXI_0_AWLOCK, // @[:@48700.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@48700.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@48700.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@48700.4]
  output         io_M_AXI_0_AWVALID, // @[:@48700.4]
  input          io_M_AXI_0_AWREADY, // @[:@48700.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@48700.4]
  output [39:0]  io_M_AXI_0_ARUSER, // @[:@48700.4]
  output [39:0]  io_M_AXI_0_ARADDR, // @[:@48700.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@48700.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@48700.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@48700.4]
  output         io_M_AXI_0_ARLOCK, // @[:@48700.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@48700.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@48700.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@48700.4]
  output         io_M_AXI_0_ARVALID, // @[:@48700.4]
  input          io_M_AXI_0_ARREADY, // @[:@48700.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@48700.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@48700.4]
  output         io_M_AXI_0_WLAST, // @[:@48700.4]
  output         io_M_AXI_0_WVALID, // @[:@48700.4]
  input          io_M_AXI_0_WREADY, // @[:@48700.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@48700.4]
  input  [39:0]  io_M_AXI_0_RUSER, // @[:@48700.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@48700.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@48700.4]
  input          io_M_AXI_0_RLAST, // @[:@48700.4]
  input          io_M_AXI_0_RVALID, // @[:@48700.4]
  output         io_M_AXI_0_RREADY, // @[:@48700.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@48700.4]
  input  [39:0]  io_M_AXI_0_BUSER, // @[:@48700.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@48700.4]
  input          io_M_AXI_0_BVALID, // @[:@48700.4]
  output         io_M_AXI_0_BREADY, // @[:@48700.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@48700.4]
  output [39:0]  io_M_AXI_1_AWUSER, // @[:@48700.4]
  output [39:0]  io_M_AXI_1_AWADDR, // @[:@48700.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@48700.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@48700.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@48700.4]
  output         io_M_AXI_1_AWLOCK, // @[:@48700.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@48700.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@48700.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@48700.4]
  output         io_M_AXI_1_AWVALID, // @[:@48700.4]
  input          io_M_AXI_1_AWREADY, // @[:@48700.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@48700.4]
  output [39:0]  io_M_AXI_1_ARUSER, // @[:@48700.4]
  output [39:0]  io_M_AXI_1_ARADDR, // @[:@48700.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@48700.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@48700.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@48700.4]
  output         io_M_AXI_1_ARLOCK, // @[:@48700.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@48700.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@48700.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@48700.4]
  output         io_M_AXI_1_ARVALID, // @[:@48700.4]
  input          io_M_AXI_1_ARREADY, // @[:@48700.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@48700.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@48700.4]
  output         io_M_AXI_1_WLAST, // @[:@48700.4]
  output         io_M_AXI_1_WVALID, // @[:@48700.4]
  input          io_M_AXI_1_WREADY, // @[:@48700.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@48700.4]
  input  [39:0]  io_M_AXI_1_RUSER, // @[:@48700.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@48700.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@48700.4]
  input          io_M_AXI_1_RLAST, // @[:@48700.4]
  input          io_M_AXI_1_RVALID, // @[:@48700.4]
  output         io_M_AXI_1_RREADY, // @[:@48700.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@48700.4]
  input  [39:0]  io_M_AXI_1_BUSER, // @[:@48700.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@48700.4]
  input          io_M_AXI_1_BVALID, // @[:@48700.4]
  output         io_M_AXI_1_BREADY // @[:@48700.4]
);
  wire  accel_clock; // @[Instantiator.scala 54:38:@48702.4]
  wire  accel_reset; // @[Instantiator.scala 54:38:@48702.4]
  wire  accel_io_enable; // @[Instantiator.scala 54:38:@48702.4]
  wire  accel_io_done; // @[Instantiator.scala 54:38:@48702.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 54:38:@48702.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 54:38:@48702.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 54:38:@48702.4]
  wire  FringeZynq_clock; // @[KCU1500.scala 21:24:@48792.4]
  wire  FringeZynq_reset; // @[KCU1500.scala 21:24:@48792.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 21:24:@48792.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 21:24:@48792.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[KCU1500.scala 21:24:@48792.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[KCU1500.scala 21:24:@48792.4]
  wire  FringeZynq_io_enable; // @[KCU1500.scala 21:24:@48792.4]
  wire  FringeZynq_io_done; // @[KCU1500.scala 21:24:@48792.4]
  wire  FringeZynq_io_reset; // @[KCU1500.scala 21:24:@48792.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[KCU1500.scala 21:24:@48792.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[KCU1500.scala 21:24:@48792.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[KCU1500.scala 21:24:@48792.4]
  AccelTop accel ( // @[Instantiator.scala 54:38:@48702.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits)
  );
  FringeZynq FringeZynq ( // @[KCU1500.scala 21:24:@48792.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = 1'h0; // @[KCU1500.scala 24:21:@48810.4]
  assign io_S_AXI_ARREADY = 1'h0; // @[KCU1500.scala 24:21:@48806.4]
  assign io_S_AXI_WREADY = 1'h0; // @[KCU1500.scala 24:21:@48802.4]
  assign io_S_AXI_RDATA = 64'h0; // @[KCU1500.scala 24:21:@48801.4]
  assign io_S_AXI_RRESP = 2'h0; // @[KCU1500.scala 24:21:@48800.4]
  assign io_S_AXI_RVALID = 1'h0; // @[KCU1500.scala 24:21:@48799.4]
  assign io_S_AXI_BRESP = 2'h0; // @[KCU1500.scala 24:21:@48797.4]
  assign io_S_AXI_BVALID = 1'h0; // @[KCU1500.scala 24:21:@48796.4]
  assign io_M_AXI_0_AWID = 32'h0; // @[KCU1500.scala 27:14:@48854.4]
  assign io_M_AXI_0_AWUSER = 40'h0; // @[KCU1500.scala 27:14:@48853.4]
  assign io_M_AXI_0_AWADDR = 40'h0; // @[KCU1500.scala 27:14:@48852.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[KCU1500.scala 27:14:@48851.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[KCU1500.scala 27:14:@48850.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[KCU1500.scala 27:14:@48849.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[KCU1500.scala 27:14:@48848.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[KCU1500.scala 27:14:@48847.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[KCU1500.scala 27:14:@48846.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[KCU1500.scala 27:14:@48845.4]
  assign io_M_AXI_0_AWVALID = 1'h0; // @[KCU1500.scala 27:14:@48844.4]
  assign io_M_AXI_0_ARID = 32'h0; // @[KCU1500.scala 27:14:@48842.4]
  assign io_M_AXI_0_ARUSER = 40'h0; // @[KCU1500.scala 27:14:@48841.4]
  assign io_M_AXI_0_ARADDR = 40'h0; // @[KCU1500.scala 27:14:@48840.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[KCU1500.scala 27:14:@48839.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[KCU1500.scala 27:14:@48838.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[KCU1500.scala 27:14:@48837.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[KCU1500.scala 27:14:@48836.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[KCU1500.scala 27:14:@48835.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[KCU1500.scala 27:14:@48834.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[KCU1500.scala 27:14:@48833.4]
  assign io_M_AXI_0_ARVALID = 1'h0; // @[KCU1500.scala 27:14:@48832.4]
  assign io_M_AXI_0_WDATA = 512'h0; // @[KCU1500.scala 27:14:@48830.4]
  assign io_M_AXI_0_WSTRB = 64'h0; // @[KCU1500.scala 27:14:@48829.4]
  assign io_M_AXI_0_WLAST = 1'h0; // @[KCU1500.scala 27:14:@48828.4]
  assign io_M_AXI_0_WVALID = 1'h0; // @[KCU1500.scala 27:14:@48827.4]
  assign io_M_AXI_0_RREADY = 1'h0; // @[KCU1500.scala 27:14:@48819.4]
  assign io_M_AXI_0_BREADY = 1'h0; // @[KCU1500.scala 27:14:@48814.4]
  assign io_M_AXI_1_AWID = 32'h0; // @[KCU1500.scala 27:14:@48895.4]
  assign io_M_AXI_1_AWUSER = 40'h0; // @[KCU1500.scala 27:14:@48894.4]
  assign io_M_AXI_1_AWADDR = 40'h0; // @[KCU1500.scala 27:14:@48893.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[KCU1500.scala 27:14:@48892.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[KCU1500.scala 27:14:@48891.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[KCU1500.scala 27:14:@48890.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[KCU1500.scala 27:14:@48889.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[KCU1500.scala 27:14:@48888.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[KCU1500.scala 27:14:@48887.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[KCU1500.scala 27:14:@48886.4]
  assign io_M_AXI_1_AWVALID = 1'h0; // @[KCU1500.scala 27:14:@48885.4]
  assign io_M_AXI_1_ARID = 32'h0; // @[KCU1500.scala 27:14:@48883.4]
  assign io_M_AXI_1_ARUSER = 40'h0; // @[KCU1500.scala 27:14:@48882.4]
  assign io_M_AXI_1_ARADDR = 40'h0; // @[KCU1500.scala 27:14:@48881.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[KCU1500.scala 27:14:@48880.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[KCU1500.scala 27:14:@48879.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[KCU1500.scala 27:14:@48878.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[KCU1500.scala 27:14:@48877.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[KCU1500.scala 27:14:@48876.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[KCU1500.scala 27:14:@48875.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[KCU1500.scala 27:14:@48874.4]
  assign io_M_AXI_1_ARVALID = 1'h0; // @[KCU1500.scala 27:14:@48873.4]
  assign io_M_AXI_1_WDATA = 512'h0; // @[KCU1500.scala 27:14:@48871.4]
  assign io_M_AXI_1_WSTRB = 64'h0; // @[KCU1500.scala 27:14:@48870.4]
  assign io_M_AXI_1_WLAST = 1'h0; // @[KCU1500.scala 27:14:@48869.4]
  assign io_M_AXI_1_WVALID = 1'h0; // @[KCU1500.scala 27:14:@48868.4]
  assign io_M_AXI_1_RREADY = 1'h0; // @[KCU1500.scala 27:14:@48860.4]
  assign io_M_AXI_1_BREADY = 1'h0; // @[KCU1500.scala 27:14:@48855.4]
  assign accel_clock = clock; // @[:@48703.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@48704.4 KCU1500.scala 57:17:@49150.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[KCU1500.scala 54:21:@49145.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[KCU1500.scala 37:21:@49061.4]
  assign FringeZynq_clock = clock; // @[:@48793.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@48794.4 KCU1500.scala 56:18:@49149.4]
  assign FringeZynq_io_done = accel_io_done; // @[KCU1500.scala 55:20:@49146.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[KCU1500.scala 40:26:@49063.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[KCU1500.scala 39:25:@49062.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule

